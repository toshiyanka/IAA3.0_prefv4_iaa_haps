### Tool : gds2def
### Version 14.1     Linux64
### Vendor : Apache Design, Inc. A Subsidiary of ANSYS, Inc. 
### Date : Jun 19 2014 02:20:56 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
MACRO c73p1rfshdxrom2048x16hb4img100_APACHECELL
 CLASS BLOCK ;
 ORIGIN 0 0 ;
 SIZE 75.432 BY 29.526 ;
 PIN iar[10]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 10.932 0.308 10.964 ;
 END
 END iar[10]
 PIN iar[0]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 11.674 0.308 11.706 ;
 END
 END iar[0]
 PIN iar[1]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 12.472 0.308 12.504 ;
 END
 END iar[1]
 PIN iar[2]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 13.088 0.308 13.12 ;
 END
 END iar[2]
 PIN iar[4]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 13.774 0.308 13.806 ;
 END
 END iar[4]
 PIN iar[3]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 14.404 0.308 14.436 ;
 END
 END iar[3]
 PIN iar[7]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 15.72 0.308 15.752 ;
 END
 END iar[7]
 PIN iar[6]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 16.406 0.308 16.438 ;
 END
 END iar[6]
 PIN iar[5]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 16.966 0.308 16.998 ;
 END
 END iar[5]
 PIN iar[9]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 17.764 0.308 17.796 ;
 END
 END iar[9]
 PIN iar[8]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 18.282 0.308 18.314 ;
 END
 END iar[8]
 PIN iren
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 15.146 0.308 15.178 ;
 END
 END iren
 PIN ickr
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 14.922 0.308 14.954 ;
 END
 END ickr
 PIN ipwreninb
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 28.544 0.308 28.576 ;
 END
 END ipwreninb
 PIN opwrenoutb
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 0.726 0.308 0.758 ;
 END
 END opwrenoutb
 PIN odout[0]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 0.95 0.308 0.982 ;
 END
 END odout[0]
 PIN odout[1]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 2.21 0.308 2.242 ;
 END
 END odout[1]
 PIN odout[2]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 3.456 0.308 3.488 ;
 END
 END odout[2]
 PIN odout[3]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 4.716 0.308 4.748 ;
 END
 END odout[3]
 PIN odout[4]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 5.85 0.308 5.882 ;
 END
 END odout[4]
 PIN odout[5]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 7.222 0.308 7.254 ;
 END
 END odout[5]
 PIN odout[6]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 8.482 0.308 8.514 ;
 END
 END odout[6]
 PIN odout[7]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 9.728 0.308 9.76 ;
 END
 END odout[7]
 PIN odout[8]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 19.08 0.308 19.112 ;
 END
 END odout[8]
 PIN odout[9]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 20.452 0.308 20.484 ;
 END
 END odout[9]
 PIN odout[10]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 21.698 0.308 21.73 ;
 END
 END odout[10]
 PIN odout[11]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 22.846 0.308 22.878 ;
 END
 END odout[11]
 PIN odout[12]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 24.092 0.308 24.124 ;
 END
 END odout[12]
 PIN odout[13]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 25.352 0.308 25.384 ;
 END
 END odout[13]
 PIN odout[14]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 26.836 0.308 26.868 ;
 END
 END odout[14]
 PIN odout[15]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 28.194 0.308 28.226 ;
 END
 END odout[15]
 PIN vccd_1p0
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 2.978 0.43 3.178 ;
 END
 END vccd_1p0
 PIN vccd_1p0.gds1
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 1.022 5.202 1.222 ;
 END
 END vccd_1p0.gds1
 PIN vccd_1p0.gds2
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 1.013 1.542 1.213 ;
 END
 END vccd_1p0.gds2
 PIN vccd_1p0.gds3
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 4.793 1.542 4.993 ;
 END
 END vccd_1p0.gds3
 PIN vccd_1p0.gds4
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 4.6755 5.202 4.8755 ;
 END
 END vccd_1p0.gds4
 PIN vccd_1p0.gds5
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 3.533 1.542 3.733 ;
 END
 END vccd_1p0.gds5
 PIN vccd_1p0.gds6
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 3.4155 5.202 3.6155 ;
 END
 END vccd_1p0.gds6
 PIN vccd_1p0.gds7
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 3.089 0.548 3.289 ;
 END
 END vccd_1p0.gds7
 PIN vccd_1p0.gds8
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 3.0505 0.858 3.2505 ;
 END
 END vccd_1p0.gds8
 PIN vccd_1p0.gds9
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 2.888 1.362 3.088 ;
 END
 END vccd_1p0.gds9
 PIN vccd_1p0.gds10
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 3.022 1.782 3.222 ;
 END
 END vccd_1p0.gds10
 PIN vccd_1p0.gds11
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 2.273 1.542 2.473 ;
 END
 END vccd_1p0.gds11
 PIN vccd_1p0.gds12
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 2.987 1.218 3.187 ;
 END
 END vccd_1p0.gds12
 PIN vccd_1p0.gds13
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 2.1555 5.202 2.3555 ;
 END
 END vccd_1p0.gds13
 PIN vccd_1p0.gds14
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 3.157 1.962 3.357 ;
 END
 END vccd_1p0.gds14
 PIN vccd_1p0.gds15
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 2.9685 2.202 3.1685 ;
 END
 END vccd_1p0.gds15
 PIN vccd_1p0.gds16
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 3.0145 2.462 3.2145 ;
 END
 END vccd_1p0.gds16
 PIN vccd_1p0.gds17
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 3.007 2.622 3.207 ;
 END
 END vccd_1p0.gds17
 PIN vccd_1p0.gds18
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 3.007 1.09 3.207 ;
 END
 END vccd_1p0.gds18
 PIN vccd_1p0.gds19
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 2.8915 3.042 3.0915 ;
 END
 END vccd_1p0.gds19
 PIN vccd_1p0.gds20
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 3.02 2.882 3.22 ;
 END
 END vccd_1p0.gds20
 PIN vccd_1p0.gds21
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 3.016 3.262 3.216 ;
 END
 END vccd_1p0.gds21
 PIN vccd_1p0.gds22
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 3.0585 4.738 3.2585 ;
 END
 END vccd_1p0.gds22
 PIN vccd_1p0.gds23
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 2.98 3.39 3.18 ;
 END
 END vccd_1p0.gds23
 PIN vccd_1p0.gds24
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 3.059 3.666 3.259 ;
 END
 END vccd_1p0.gds24
 PIN vccd_1p0.gds25
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 3.0725 4.066 3.2725 ;
 END
 END vccd_1p0.gds25
 PIN vccd_1p0.gds26
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 3.0725 3.858 3.2725 ;
 END
 END vccd_1p0.gds26
 PIN vccd_1p0.gds27
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 3.058 4.546 3.258 ;
 END
 END vccd_1p0.gds27
 PIN vccd_1p0.gds28
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 3.02 4.258 3.22 ;
 END
 END vccd_1p0.gds28
 PIN vccd_1p0.gds29
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 3.082 5.01 3.282 ;
 END
 END vccd_1p0.gds29
 PIN vccd_1p0.gds30
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 3.584 1.0395 3.64 1.2395 ;
 RECT 3.584 2.2995 3.64 2.4995 ;
 RECT 3.584 3.5595 3.64 3.7595 ;
 RECT 3.584 4.8195 3.64 5.0195 ;
 RECT 4.34 4.918 4.396 5.118 ;
 RECT 4.172 4.918 4.228 5.118 ;
 RECT 4.76 4.8775 4.816 5.0775 ;
 RECT 5.096 4.918 5.152 5.118 ;
 RECT 4.928 4.8775 4.984 5.0775 ;
 RECT 4.34 3.658 4.396 3.858 ;
 RECT 4.172 3.658 4.228 3.858 ;
 RECT 4.76 3.6175 4.816 3.8175 ;
 RECT 5.096 3.658 5.152 3.858 ;
 RECT 4.928 3.6175 4.984 3.8175 ;
 RECT 4.34 2.398 4.396 2.598 ;
 RECT 4.172 2.398 4.228 2.598 ;
 RECT 4.76 2.3575 4.816 2.5575 ;
 RECT 5.096 2.398 5.152 2.598 ;
 RECT 4.928 2.3575 4.984 2.5575 ;
 RECT 4.34 1.138 4.396 1.338 ;
 RECT 4.172 1.138 4.228 1.338 ;
 RECT 4.76 1.0975 4.816 1.2975 ;
 RECT 5.096 1.138 5.152 1.338 ;
 RECT 4.928 1.0975 4.984 1.2975 ;
 END
 END vccd_1p0.gds30
 PIN vccd_1p0.gds31
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 3.0725 6.838 3.2725 ;
 END
 END vccd_1p0.gds31
 PIN vccd_1p0.gds32
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 3.082 6.05 3.282 ;
 END
 END vccd_1p0.gds32
 PIN vccd_1p0.gds33
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.754 3.02 5.794 3.22 ;
 END
 END vccd_1p0.gds33
 PIN vccd_1p0.gds34
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 3.109 6.306 3.309 ;
 END
 END vccd_1p0.gds34
 PIN vccd_1p0.gds35
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 3.0725 5.41 3.2725 ;
 END
 END vccd_1p0.gds35
 PIN vccd_1p0.gds36
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 3.0725 5.922 3.2725 ;
 END
 END vccd_1p0.gds36
 PIN vccd_1p0.gds37
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 2.962 5.602 3.162 ;
 END
 END vccd_1p0.gds37
 PIN vccd_1p0.gds38
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 2.999 6.582 3.199 ;
 END
 END vccd_1p0.gds38
 PIN vccd_1p0.gds39
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.6 4.918 5.656 5.118 ;
 RECT 5.432 4.8295 5.488 5.0295 ;
 RECT 5.264 4.918 5.32 5.118 ;
 RECT 5.936 4.8295 5.992 5.0295 ;
 RECT 5.768 4.8295 5.824 5.0295 ;
 RECT 6.44 4.8465 6.496 5.0465 ;
 RECT 6.272 4.8295 6.328 5.0295 ;
 RECT 6.104 4.918 6.16 5.118 ;
 RECT 5.6 3.658 5.656 3.858 ;
 RECT 5.432 3.5695 5.488 3.7695 ;
 RECT 5.264 3.658 5.32 3.858 ;
 RECT 5.936 3.5695 5.992 3.7695 ;
 RECT 5.768 3.5695 5.824 3.7695 ;
 RECT 6.44 3.5865 6.496 3.7865 ;
 RECT 6.272 3.5695 6.328 3.7695 ;
 RECT 6.104 3.658 6.16 3.858 ;
 RECT 5.6 2.398 5.656 2.598 ;
 RECT 5.432 2.3095 5.488 2.5095 ;
 RECT 5.264 2.398 5.32 2.598 ;
 RECT 5.936 2.3095 5.992 2.5095 ;
 RECT 5.768 2.3095 5.824 2.5095 ;
 RECT 6.44 2.3265 6.496 2.5265 ;
 RECT 6.272 2.3095 6.328 2.5095 ;
 RECT 6.104 2.398 6.16 2.598 ;
 RECT 5.6 1.138 5.656 1.338 ;
 RECT 5.432 1.0495 5.488 1.2495 ;
 RECT 5.264 1.138 5.32 1.338 ;
 RECT 5.936 1.0495 5.992 1.2495 ;
 RECT 5.768 1.0495 5.824 1.2495 ;
 RECT 6.44 1.0665 6.496 1.2665 ;
 RECT 6.272 1.0495 6.328 1.2495 ;
 RECT 6.104 1.138 6.16 1.338 ;
 END
 END vccd_1p0.gds39
 PIN vccd_1p0.gds40
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 1.36 13.978 1.56 ;
 END
 END vccd_1p0.gds40
 PIN vccd_1p0.gds41
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 2.62 13.978 2.82 ;
 END
 END vccd_1p0.gds41
 PIN vccd_1p0.gds42
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 3.88 13.978 4.08 ;
 END
 END vccd_1p0.gds42
 PIN vccd_1p0.gds43
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 1.36 14.398 1.56 ;
 END
 END vccd_1p0.gds43
 PIN vccd_1p0.gds44
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 2.62 14.398 2.82 ;
 END
 END vccd_1p0.gds44
 PIN vccd_1p0.gds45
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 5.14 13.978 5.34 ;
 END
 END vccd_1p0.gds45
 PIN vccd_1p0.gds46
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 5.14 14.398 5.34 ;
 END
 END vccd_1p0.gds46
 PIN vccd_1p0.gds47
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 5.2675 14.934 5.4675 ;
 END
 END vccd_1p0.gds47
 PIN vccd_1p0.gds48
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 2.82 13.738 3.02 ;
 END
 END vccd_1p0.gds48
 PIN vccd_1p0.gds49
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 2.8975 13.138 3.0975 ;
 END
 END vccd_1p0.gds49
 PIN vccd_1p0.gds50
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 3.88 14.398 4.08 ;
 END
 END vccd_1p0.gds50
 PIN vccd_1p0.gds51
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 4.0075 14.934 4.2075 ;
 END
 END vccd_1p0.gds51
 PIN vccd_1p0.gds52
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 3.072 14.742 3.272 ;
 END
 END vccd_1p0.gds52
 PIN vccd_1p0.gds53
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 3.02 12.898 3.22 ;
 END
 END vccd_1p0.gds53
 PIN vccd_1p0.gds54
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 3.016 12.654 3.216 ;
 END
 END vccd_1p0.gds54
 PIN vccd_1p0.gds55
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 2.9745 12.526 3.1745 ;
 END
 END vccd_1p0.gds55
 PIN vccd_1p0.gds56
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 2.7475 14.934 2.9475 ;
 END
 END vccd_1p0.gds56
 PIN vccd_1p0.gds57
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 1.4875 14.934 1.6875 ;
 END
 END vccd_1p0.gds57
 PIN vccd_1p0.gds58
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 1.424 16.226 1.624 ;
 END
 END vccd_1p0.gds58
 PIN vccd_1p0.gds59
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 2.684 16.226 2.884 ;
 END
 END vccd_1p0.gds59
 PIN vccd_1p0.gds60
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 3.944 16.226 4.144 ;
 END
 END vccd_1p0.gds60
 PIN vccd_1p0.gds61
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 5.204 16.226 5.404 ;
 END
 END vccd_1p0.gds61
 PIN vccd_1p0.gds62
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 3.072 15.29 3.272 ;
 END
 END vccd_1p0.gds62
 PIN vccd_1p0.gds63
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 2.9985 17.574 3.1985 ;
 END
 END vccd_1p0.gds63
 PIN vccd_1p0.gds64
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 3.054 15.742 3.254 ;
 END
 END vccd_1p0.gds64
 PIN vccd_1p0.gds65
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 3.054 15.498 3.254 ;
 END
 END vccd_1p0.gds65
 PIN vccd_1p0.gds66
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 3.02 17.734 3.22 ;
 END
 END vccd_1p0.gds66
 PIN vccd_1p0.gds67
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 2.9235 17.154 3.1235 ;
 END
 END vccd_1p0.gds67
 PIN vccd_1p0.gds68
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 2.9745 18.09 3.1745 ;
 END
 END vccd_1p0.gds68
 PIN vccd_1p0.gds69
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 3.016 17.962 3.216 ;
 END
 END vccd_1p0.gds69
 PIN vccd_1p0.gds70
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 2.9785 23.842 3.1785 ;
 END
 END vccd_1p0.gds70
 PIN vccd_1p0.gds71
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 3.02 29.95 3.22 ;
 END
 END vccd_1p0.gds71
 PIN vccd_1p0.gds72
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 3.016 29.706 3.216 ;
 END
 END vccd_1p0.gds72
 PIN vccd_1p0.gds73
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 2.9745 29.578 3.1745 ;
 END
 END vccd_1p0.gds73
 PIN vccd_1p0.gds74
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 1.36 31.03 1.56 ;
 END
 END vccd_1p0.gds74
 PIN vccd_1p0.gds75
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 2.62 31.03 2.82 ;
 END
 END vccd_1p0.gds75
 PIN vccd_1p0.gds76
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 3.88 31.03 4.08 ;
 END
 END vccd_1p0.gds76
 PIN vccd_1p0.gds77
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 5.14 31.03 5.34 ;
 END
 END vccd_1p0.gds77
 PIN vccd_1p0.gds78
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 1.424 33.278 1.624 ;
 END
 END vccd_1p0.gds78
 PIN vccd_1p0.gds79
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 5.204 33.278 5.404 ;
 END
 END vccd_1p0.gds79
 PIN vccd_1p0.gds80
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 5.14 31.45 5.34 ;
 END
 END vccd_1p0.gds80
 PIN vccd_1p0.gds81
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 5.2675 31.986 5.4675 ;
 END
 END vccd_1p0.gds81
 PIN vccd_1p0.gds82
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 3.944 33.278 4.144 ;
 END
 END vccd_1p0.gds82
 PIN vccd_1p0.gds83
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 3.88 31.45 4.08 ;
 END
 END vccd_1p0.gds83
 PIN vccd_1p0.gds84
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 4.0075 31.986 4.2075 ;
 END
 END vccd_1p0.gds84
 PIN vccd_1p0.gds85
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 2.684 33.278 2.884 ;
 END
 END vccd_1p0.gds85
 PIN vccd_1p0.gds86
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 2.62 31.45 2.82 ;
 END
 END vccd_1p0.gds86
 PIN vccd_1p0.gds87
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 2.7475 31.986 2.9475 ;
 END
 END vccd_1p0.gds87
 PIN vccd_1p0.gds88
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 3.054 32.794 3.254 ;
 END
 END vccd_1p0.gds88
 PIN vccd_1p0.gds89
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 3.072 32.342 3.272 ;
 END
 END vccd_1p0.gds89
 PIN vccd_1p0.gds90
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 1.36 31.45 1.56 ;
 END
 END vccd_1p0.gds90
 PIN vccd_1p0.gds91
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 1.4875 31.986 1.6875 ;
 END
 END vccd_1p0.gds91
 PIN vccd_1p0.gds92
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 3.072 31.794 3.272 ;
 END
 END vccd_1p0.gds92
 PIN vccd_1p0.gds93
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 2.953 34.626 3.153 ;
 END
 END vccd_1p0.gds93
 PIN vccd_1p0.gds94
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 2.9745 35.142 3.1745 ;
 END
 END vccd_1p0.gds94
 PIN vccd_1p0.gds95
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 3.016 35.014 3.216 ;
 END
 END vccd_1p0.gds95
 PIN vccd_1p0.gds96
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 2.82 30.79 3.02 ;
 END
 END vccd_1p0.gds96
 PIN vccd_1p0.gds97
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 2.8975 30.19 3.0975 ;
 END
 END vccd_1p0.gds97
 PIN vccd_1p0.gds98
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 2.9235 34.206 3.1235 ;
 END
 END vccd_1p0.gds98
 PIN vccd_1p0.gds99
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 3.0725 34.786 3.2725 ;
 END
 END vccd_1p0.gds99
 PIN vccd_1p0.gds100
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 3.054 32.55 3.254 ;
 END
 END vccd_1p0.gds100
 PIN vccd_1p0.gds101
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 2.9785 40.894 3.1785 ;
 END
 END vccd_1p0.gds101
 PIN vccd_1p0.gds102
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 1.36 48.082 1.56 ;
 END
 END vccd_1p0.gds102
 PIN vccd_1p0.gds103
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 2.62 48.082 2.82 ;
 END
 END vccd_1p0.gds103
 PIN vccd_1p0.gds104
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 5.14 48.082 5.34 ;
 END
 END vccd_1p0.gds104
 PIN vccd_1p0.gds105
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 3.88 48.082 4.08 ;
 END
 END vccd_1p0.gds105
 PIN vccd_1p0.gds106
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 2.82 47.842 3.02 ;
 END
 END vccd_1p0.gds106
 PIN vccd_1p0.gds107
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 2.8975 47.242 3.0975 ;
 END
 END vccd_1p0.gds107
 PIN vccd_1p0.gds108
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 1.36 48.502 1.56 ;
 END
 END vccd_1p0.gds108
 PIN vccd_1p0.gds109
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 2.62 48.502 2.82 ;
 END
 END vccd_1p0.gds109
 PIN vccd_1p0.gds110
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 5.14 48.502 5.34 ;
 END
 END vccd_1p0.gds110
 PIN vccd_1p0.gds111
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 5.2675 49.038 5.4675 ;
 END
 END vccd_1p0.gds111
 PIN vccd_1p0.gds112
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 3.072 49.394 3.272 ;
 END
 END vccd_1p0.gds112
 PIN vccd_1p0.gds113
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 3.072 48.846 3.272 ;
 END
 END vccd_1p0.gds113
 PIN vccd_1p0.gds114
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 3.88 48.502 4.08 ;
 END
 END vccd_1p0.gds114
 PIN vccd_1p0.gds115
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 4.0075 49.038 4.2075 ;
 END
 END vccd_1p0.gds115
 PIN vccd_1p0.gds116
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 2.7475 49.038 2.9475 ;
 END
 END vccd_1p0.gds116
 PIN vccd_1p0.gds117
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 3.054 49.846 3.254 ;
 END
 END vccd_1p0.gds117
 PIN vccd_1p0.gds118
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 3.054 49.602 3.254 ;
 END
 END vccd_1p0.gds118
 PIN vccd_1p0.gds119
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 1.4875 49.038 1.6875 ;
 END
 END vccd_1p0.gds119
 PIN vccd_1p0.gds120
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 3.02 47.002 3.22 ;
 END
 END vccd_1p0.gds120
 PIN vccd_1p0.gds121
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 3.016 46.758 3.216 ;
 END
 END vccd_1p0.gds121
 PIN vccd_1p0.gds122
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 2.9745 46.63 3.1745 ;
 END
 END vccd_1p0.gds122
 PIN vccd_1p0.gds123
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 1.424 50.33 1.624 ;
 END
 END vccd_1p0.gds123
 PIN vccd_1p0.gds124
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 2.684 50.33 2.884 ;
 END
 END vccd_1p0.gds124
 PIN vccd_1p0.gds125
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 3.944 50.33 4.144 ;
 END
 END vccd_1p0.gds125
 PIN vccd_1p0.gds126
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 5.204 50.33 5.404 ;
 END
 END vccd_1p0.gds126
 PIN vccd_1p0.gds127
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 2.9985 51.678 3.1985 ;
 END
 END vccd_1p0.gds127
 PIN vccd_1p0.gds128
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 2.9745 52.194 3.1745 ;
 END
 END vccd_1p0.gds128
 PIN vccd_1p0.gds129
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 3.016 52.066 3.216 ;
 END
 END vccd_1p0.gds129
 PIN vccd_1p0.gds130
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 2.9235 51.258 3.1235 ;
 END
 END vccd_1p0.gds130
 PIN vccd_1p0.gds131
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 3.02 51.838 3.22 ;
 END
 END vccd_1p0.gds131
 PIN vccd_1p0.gds132
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 2.9785 57.946 3.1785 ;
 END
 END vccd_1p0.gds132
 PIN vccd_1p0.gds133
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 1.36 65.134 1.56 ;
 END
 END vccd_1p0.gds133
 PIN vccd_1p0.gds134
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 2.62 65.134 2.82 ;
 END
 END vccd_1p0.gds134
 PIN vccd_1p0.gds135
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 3.88 65.134 4.08 ;
 END
 END vccd_1p0.gds135
 PIN vccd_1p0.gds136
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 5.14 65.134 5.34 ;
 END
 END vccd_1p0.gds136
 PIN vccd_1p0.gds137
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 2.82 64.894 3.02 ;
 END
 END vccd_1p0.gds137
 PIN vccd_1p0.gds138
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 2.8975 64.294 3.0975 ;
 END
 END vccd_1p0.gds138
 PIN vccd_1p0.gds139
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 3.02 64.054 3.22 ;
 END
 END vccd_1p0.gds139
 PIN vccd_1p0.gds140
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 3.016 63.81 3.216 ;
 END
 END vccd_1p0.gds140
 PIN vccd_1p0.gds141
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 2.9745 63.682 3.1745 ;
 END
 END vccd_1p0.gds141
 PIN vccd_1p0.gds142
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 1.424 67.382 1.624 ;
 END
 END vccd_1p0.gds142
 PIN vccd_1p0.gds143
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 1.36 65.554 1.56 ;
 END
 END vccd_1p0.gds143
 PIN vccd_1p0.gds144
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 2.684 67.382 2.884 ;
 END
 END vccd_1p0.gds144
 PIN vccd_1p0.gds145
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 2.62 65.554 2.82 ;
 END
 END vccd_1p0.gds145
 PIN vccd_1p0.gds146
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 3.944 67.382 4.144 ;
 END
 END vccd_1p0.gds146
 PIN vccd_1p0.gds147
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 5.204 67.382 5.404 ;
 END
 END vccd_1p0.gds147
 PIN vccd_1p0.gds148
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 5.14 65.554 5.34 ;
 END
 END vccd_1p0.gds148
 PIN vccd_1p0.gds149
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 5.2675 66.09 5.4675 ;
 END
 END vccd_1p0.gds149
 PIN vccd_1p0.gds150
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 3.072 66.446 3.272 ;
 END
 END vccd_1p0.gds150
 PIN vccd_1p0.gds151
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 3.072 65.898 3.272 ;
 END
 END vccd_1p0.gds151
 PIN vccd_1p0.gds152
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 3.88 65.554 4.08 ;
 END
 END vccd_1p0.gds152
 PIN vccd_1p0.gds153
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 4.0075 66.09 4.2075 ;
 END
 END vccd_1p0.gds153
 PIN vccd_1p0.gds154
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 2.9985 68.73 3.1985 ;
 END
 END vccd_1p0.gds154
 PIN vccd_1p0.gds155
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 2.9745 69.246 3.1745 ;
 END
 END vccd_1p0.gds155
 PIN vccd_1p0.gds156
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 3.016 69.118 3.216 ;
 END
 END vccd_1p0.gds156
 PIN vccd_1p0.gds157
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 2.9235 68.31 3.1235 ;
 END
 END vccd_1p0.gds157
 PIN vccd_1p0.gds158
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 2.7475 66.09 2.9475 ;
 END
 END vccd_1p0.gds158
 PIN vccd_1p0.gds159
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 3.054 66.898 3.254 ;
 END
 END vccd_1p0.gds159
 PIN vccd_1p0.gds160
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 3.054 66.654 3.254 ;
 END
 END vccd_1p0.gds160
 PIN vccd_1p0.gds161
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 1.4875 66.09 1.6875 ;
 END
 END vccd_1p0.gds161
 PIN vccd_1p0.gds162
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 3.02 68.89 3.22 ;
 END
 END vccd_1p0.gds162
 PIN vccd_1p0.gds163
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 8.018 0.43 8.218 ;
 END
 END vccd_1p0.gds163
 PIN vccd_1p0.gds164
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 7.313 1.542 7.513 ;
 END
 END vccd_1p0.gds164
 PIN vccd_1p0.gds165
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 7.1955 5.202 7.3955 ;
 END
 END vccd_1p0.gds165
 PIN vccd_1p0.gds166
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 6.053 1.542 6.253 ;
 END
 END vccd_1p0.gds166
 PIN vccd_1p0.gds167
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 5.9355 5.202 6.1355 ;
 END
 END vccd_1p0.gds167
 PIN vccd_1p0.gds168
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 8.573 1.542 8.773 ;
 END
 END vccd_1p0.gds168
 PIN vccd_1p0.gds169
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 8.4555 5.202 8.6555 ;
 END
 END vccd_1p0.gds169
 PIN vccd_1p0.gds170
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 8.414 0.548 8.614 ;
 END
 END vccd_1p0.gds170
 PIN vccd_1p0.gds171
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 8.0905 0.858 8.2905 ;
 END
 END vccd_1p0.gds171
 PIN vccd_1p0.gds172
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 7.928 1.362 8.128 ;
 END
 END vccd_1p0.gds172
 PIN vccd_1p0.gds173
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 8.13 1.782 8.33 ;
 END
 END vccd_1p0.gds173
 PIN vccd_1p0.gds174
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 8.027 1.218 8.227 ;
 END
 END vccd_1p0.gds174
 PIN vccd_1p0.gds175
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 9.833 1.542 10.033 ;
 END
 END vccd_1p0.gds175
 PIN vccd_1p0.gds176
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 8.2955 1.962 8.4955 ;
 END
 END vccd_1p0.gds176
 PIN vccd_1p0.gds177
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 8.0085 2.202 8.2085 ;
 END
 END vccd_1p0.gds177
 PIN vccd_1p0.gds178
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 8.0545 2.462 8.2545 ;
 END
 END vccd_1p0.gds178
 PIN vccd_1p0.gds179
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 8.047 2.622 8.247 ;
 END
 END vccd_1p0.gds179
 PIN vccd_1p0.gds180
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 8.047 1.09 8.247 ;
 END
 END vccd_1p0.gds180
 PIN vccd_1p0.gds181
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 7.9315 3.042 8.1315 ;
 END
 END vccd_1p0.gds181
 PIN vccd_1p0.gds182
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 8.06 2.882 8.26 ;
 END
 END vccd_1p0.gds182
 PIN vccd_1p0.gds183
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 8.056 3.262 8.256 ;
 END
 END vccd_1p0.gds183
 PIN vccd_1p0.gds184
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 8.0985 4.738 8.2985 ;
 END
 END vccd_1p0.gds184
 PIN vccd_1p0.gds185
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 9.805 5.202 10.005 ;
 END
 END vccd_1p0.gds185
 PIN vccd_1p0.gds186
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 8.02 3.39 8.22 ;
 END
 END vccd_1p0.gds186
 PIN vccd_1p0.gds187
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 8.099 3.666 8.299 ;
 END
 END vccd_1p0.gds187
 PIN vccd_1p0.gds188
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 8.1125 4.066 8.3125 ;
 END
 END vccd_1p0.gds188
 PIN vccd_1p0.gds189
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 8.1125 3.858 8.3125 ;
 END
 END vccd_1p0.gds189
 PIN vccd_1p0.gds190
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 8.165 4.546 8.365 ;
 END
 END vccd_1p0.gds190
 PIN vccd_1p0.gds191
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 8.06 4.258 8.26 ;
 END
 END vccd_1p0.gds191
 PIN vccd_1p0.gds192
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 8.122 5.01 8.322 ;
 END
 END vccd_1p0.gds192
 PIN vccd_1p0.gds193
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 3.584 6.0795 3.64 6.2795 ;
 RECT 3.584 7.3395 3.64 7.5395 ;
 RECT 3.584 8.5995 3.64 8.7995 ;
 RECT 3.584 9.8595 3.64 10.0595 ;
 RECT 4.34 9.958 4.396 10.158 ;
 RECT 4.172 9.958 4.228 10.158 ;
 RECT 4.76 9.9175 4.816 10.1175 ;
 RECT 5.096 9.958 5.152 10.158 ;
 RECT 4.928 9.9175 4.984 10.1175 ;
 RECT 4.34 8.698 4.396 8.898 ;
 RECT 4.172 8.698 4.228 8.898 ;
 RECT 4.76 8.6575 4.816 8.8575 ;
 RECT 5.096 8.698 5.152 8.898 ;
 RECT 4.928 8.6575 4.984 8.8575 ;
 RECT 4.34 7.438 4.396 7.638 ;
 RECT 4.172 7.438 4.228 7.638 ;
 RECT 4.76 7.3975 4.816 7.5975 ;
 RECT 5.096 7.438 5.152 7.638 ;
 RECT 4.928 7.3975 4.984 7.5975 ;
 RECT 4.34 6.178 4.396 6.378 ;
 RECT 4.172 6.178 4.228 6.378 ;
 RECT 4.76 6.1375 4.816 6.3375 ;
 RECT 5.096 6.178 5.152 6.378 ;
 RECT 4.928 6.1375 4.984 6.3375 ;
 END
 END vccd_1p0.gds193
 PIN vccd_1p0.gds194
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 8.1125 6.838 8.3125 ;
 END
 END vccd_1p0.gds194
 PIN vccd_1p0.gds195
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 8.122 6.05 8.322 ;
 END
 END vccd_1p0.gds195
 PIN vccd_1p0.gds196
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.754 8.06 5.794 8.26 ;
 END
 END vccd_1p0.gds196
 PIN vccd_1p0.gds197
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 8.149 6.306 8.349 ;
 END
 END vccd_1p0.gds197
 PIN vccd_1p0.gds198
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 8.1125 5.41 8.3125 ;
 END
 END vccd_1p0.gds198
 PIN vccd_1p0.gds199
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 8.1125 5.922 8.3125 ;
 END
 END vccd_1p0.gds199
 PIN vccd_1p0.gds200
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 8.08 5.602 8.28 ;
 END
 END vccd_1p0.gds200
 PIN vccd_1p0.gds201
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 8.039 6.582 8.239 ;
 END
 END vccd_1p0.gds201
 PIN vccd_1p0.gds202
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.6 9.958 5.656 10.158 ;
 RECT 5.432 9.8695 5.488 10.0695 ;
 RECT 5.264 9.958 5.32 10.158 ;
 RECT 5.936 9.8695 5.992 10.0695 ;
 RECT 5.768 9.8695 5.824 10.0695 ;
 RECT 6.44 9.8865 6.496 10.0865 ;
 RECT 6.272 9.8695 6.328 10.0695 ;
 RECT 6.104 9.958 6.16 10.158 ;
 RECT 5.6 8.698 5.656 8.898 ;
 RECT 5.432 8.6095 5.488 8.8095 ;
 RECT 5.264 8.698 5.32 8.898 ;
 RECT 5.936 8.6095 5.992 8.8095 ;
 RECT 5.768 8.6095 5.824 8.8095 ;
 RECT 6.44 8.6265 6.496 8.8265 ;
 RECT 6.272 8.6095 6.328 8.8095 ;
 RECT 6.104 8.698 6.16 8.898 ;
 RECT 5.6 7.438 5.656 7.638 ;
 RECT 5.432 7.3495 5.488 7.5495 ;
 RECT 5.264 7.438 5.32 7.638 ;
 RECT 5.936 7.3495 5.992 7.5495 ;
 RECT 5.768 7.3495 5.824 7.5495 ;
 RECT 6.44 7.3665 6.496 7.5665 ;
 RECT 6.272 7.3495 6.328 7.5495 ;
 RECT 6.104 7.438 6.16 7.638 ;
 RECT 5.6 6.178 5.656 6.378 ;
 RECT 5.432 6.0895 5.488 6.2895 ;
 RECT 5.264 6.178 5.32 6.378 ;
 RECT 5.936 6.0895 5.992 6.2895 ;
 RECT 5.768 6.0895 5.824 6.2895 ;
 RECT 6.44 6.1065 6.496 6.3065 ;
 RECT 6.272 6.0895 6.328 6.2895 ;
 RECT 6.104 6.178 6.16 6.378 ;
 END
 END vccd_1p0.gds202
 PIN vccd_1p0.gds203
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 8.92 13.978 9.12 ;
 END
 END vccd_1p0.gds203
 PIN vccd_1p0.gds204
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 10.18 13.978 10.38 ;
 END
 END vccd_1p0.gds204
 PIN vccd_1p0.gds205
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 8.92 14.398 9.12 ;
 END
 END vccd_1p0.gds205
 PIN vccd_1p0.gds206
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 7.66 13.978 7.86 ;
 END
 END vccd_1p0.gds206
 PIN vccd_1p0.gds207
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 6.4 14.398 6.6 ;
 END
 END vccd_1p0.gds207
 PIN vccd_1p0.gds208
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 6.5275 14.934 6.7275 ;
 END
 END vccd_1p0.gds208
 PIN vccd_1p0.gds209
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 6.4 13.978 6.6 ;
 END
 END vccd_1p0.gds209
 PIN vccd_1p0.gds210
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 7.86 13.738 8.06 ;
 END
 END vccd_1p0.gds210
 PIN vccd_1p0.gds211
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 7.9375 13.138 8.1375 ;
 END
 END vccd_1p0.gds211
 PIN vccd_1p0.gds212
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 7.66 14.398 7.86 ;
 END
 END vccd_1p0.gds212
 PIN vccd_1p0.gds213
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 7.7875 14.934 7.9875 ;
 END
 END vccd_1p0.gds213
 PIN vccd_1p0.gds214
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 10.3005 14.398 10.5005 ;
 END
 END vccd_1p0.gds214
 PIN vccd_1p0.gds215
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 10.4255 14.934 10.6255 ;
 END
 END vccd_1p0.gds215
 PIN vccd_1p0.gds216
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 8.112 14.742 8.312 ;
 END
 END vccd_1p0.gds216
 PIN vccd_1p0.gds217
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 8.06 12.898 8.26 ;
 END
 END vccd_1p0.gds217
 PIN vccd_1p0.gds218
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 8.056 12.654 8.256 ;
 END
 END vccd_1p0.gds218
 PIN vccd_1p0.gds219
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 8.0145 12.526 8.2145 ;
 END
 END vccd_1p0.gds219
 PIN vccd_1p0.gds220
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 9.0475 14.934 9.2475 ;
 END
 END vccd_1p0.gds220
 PIN vccd_1p0.gds221
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 8.984 16.226 9.184 ;
 END
 END vccd_1p0.gds221
 PIN vccd_1p0.gds222
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 6.464 16.226 6.664 ;
 END
 END vccd_1p0.gds222
 PIN vccd_1p0.gds223
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 7.724 16.226 7.924 ;
 END
 END vccd_1p0.gds223
 PIN vccd_1p0.gds224
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 8.112 15.29 8.312 ;
 END
 END vccd_1p0.gds224
 PIN vccd_1p0.gds225
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 8.0385 17.574 8.2385 ;
 END
 END vccd_1p0.gds225
 PIN vccd_1p0.gds226
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 8.094 15.742 8.294 ;
 END
 END vccd_1p0.gds226
 PIN vccd_1p0.gds227
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 8.094 15.498 8.294 ;
 END
 END vccd_1p0.gds227
 PIN vccd_1p0.gds228
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 8.06 17.734 8.26 ;
 END
 END vccd_1p0.gds228
 PIN vccd_1p0.gds229
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 7.9635 17.154 8.1635 ;
 END
 END vccd_1p0.gds229
 PIN vccd_1p0.gds230
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 8.0145 18.09 8.2145 ;
 END
 END vccd_1p0.gds230
 PIN vccd_1p0.gds231
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 8.056 17.962 8.256 ;
 END
 END vccd_1p0.gds231
 PIN vccd_1p0.gds232
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 8.0185 23.842 8.2185 ;
 END
 END vccd_1p0.gds232
 PIN vccd_1p0.gds233
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 8.06 29.95 8.26 ;
 END
 END vccd_1p0.gds233
 PIN vccd_1p0.gds234
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 8.056 29.706 8.256 ;
 END
 END vccd_1p0.gds234
 PIN vccd_1p0.gds235
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 8.0145 29.578 8.2145 ;
 END
 END vccd_1p0.gds235
 PIN vccd_1p0.gds236
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 8.92 31.03 9.12 ;
 END
 END vccd_1p0.gds236
 PIN vccd_1p0.gds237
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 10.18 31.03 10.38 ;
 END
 END vccd_1p0.gds237
 PIN vccd_1p0.gds238
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 6.4 31.03 6.6 ;
 END
 END vccd_1p0.gds238
 PIN vccd_1p0.gds239
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 8.984 33.278 9.184 ;
 END
 END vccd_1p0.gds239
 PIN vccd_1p0.gds240
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 8.92 31.45 9.12 ;
 END
 END vccd_1p0.gds240
 PIN vccd_1p0.gds241
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 7.724 33.278 7.924 ;
 END
 END vccd_1p0.gds241
 PIN vccd_1p0.gds242
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 6.464 33.278 6.664 ;
 END
 END vccd_1p0.gds242
 PIN vccd_1p0.gds243
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 6.4 31.45 6.6 ;
 END
 END vccd_1p0.gds243
 PIN vccd_1p0.gds244
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 6.5275 31.986 6.7275 ;
 END
 END vccd_1p0.gds244
 PIN vccd_1p0.gds245
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 8.094 32.794 8.294 ;
 END
 END vccd_1p0.gds245
 PIN vccd_1p0.gds246
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 7.66 31.45 7.86 ;
 END
 END vccd_1p0.gds246
 PIN vccd_1p0.gds247
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 7.7875 31.986 7.9875 ;
 END
 END vccd_1p0.gds247
 PIN vccd_1p0.gds248
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 8.112 32.342 8.312 ;
 END
 END vccd_1p0.gds248
 PIN vccd_1p0.gds249
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 8.112 31.794 8.312 ;
 END
 END vccd_1p0.gds249
 PIN vccd_1p0.gds250
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 10.3005 31.45 10.5005 ;
 END
 END vccd_1p0.gds250
 PIN vccd_1p0.gds251
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 10.4255 31.986 10.6255 ;
 END
 END vccd_1p0.gds251
 PIN vccd_1p0.gds252
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 7.993 34.626 8.193 ;
 END
 END vccd_1p0.gds252
 PIN vccd_1p0.gds253
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 9.0475 31.986 9.2475 ;
 END
 END vccd_1p0.gds253
 PIN vccd_1p0.gds254
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 8.0145 35.142 8.2145 ;
 END
 END vccd_1p0.gds254
 PIN vccd_1p0.gds255
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 8.056 35.014 8.256 ;
 END
 END vccd_1p0.gds255
 PIN vccd_1p0.gds256
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 7.66 31.03 7.86 ;
 END
 END vccd_1p0.gds256
 PIN vccd_1p0.gds257
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 7.86 30.79 8.06 ;
 END
 END vccd_1p0.gds257
 PIN vccd_1p0.gds258
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 7.9375 30.19 8.1375 ;
 END
 END vccd_1p0.gds258
 PIN vccd_1p0.gds259
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 7.9635 34.206 8.1635 ;
 END
 END vccd_1p0.gds259
 PIN vccd_1p0.gds260
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 8.1125 34.786 8.3125 ;
 END
 END vccd_1p0.gds260
 PIN vccd_1p0.gds261
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 8.094 32.55 8.294 ;
 END
 END vccd_1p0.gds261
 PIN vccd_1p0.gds262
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 8.0185 40.894 8.2185 ;
 END
 END vccd_1p0.gds262
 PIN vccd_1p0.gds263
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 8.92 48.082 9.12 ;
 END
 END vccd_1p0.gds263
 PIN vccd_1p0.gds264
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 10.18 48.082 10.38 ;
 END
 END vccd_1p0.gds264
 PIN vccd_1p0.gds265
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 7.66 48.082 7.86 ;
 END
 END vccd_1p0.gds265
 PIN vccd_1p0.gds266
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 6.4 48.082 6.6 ;
 END
 END vccd_1p0.gds266
 PIN vccd_1p0.gds267
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 7.86 47.842 8.06 ;
 END
 END vccd_1p0.gds267
 PIN vccd_1p0.gds268
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 7.9375 47.242 8.1375 ;
 END
 END vccd_1p0.gds268
 PIN vccd_1p0.gds269
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 8.92 48.502 9.12 ;
 END
 END vccd_1p0.gds269
 PIN vccd_1p0.gds270
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 7.66 48.502 7.86 ;
 END
 END vccd_1p0.gds270
 PIN vccd_1p0.gds271
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 7.7875 49.038 7.9875 ;
 END
 END vccd_1p0.gds271
 PIN vccd_1p0.gds272
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 6.4 48.502 6.6 ;
 END
 END vccd_1p0.gds272
 PIN vccd_1p0.gds273
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 6.5275 49.038 6.7275 ;
 END
 END vccd_1p0.gds273
 PIN vccd_1p0.gds274
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 8.112 49.394 8.312 ;
 END
 END vccd_1p0.gds274
 PIN vccd_1p0.gds275
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 10.3005 48.502 10.5005 ;
 END
 END vccd_1p0.gds275
 PIN vccd_1p0.gds276
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 10.4255 49.038 10.6255 ;
 END
 END vccd_1p0.gds276
 PIN vccd_1p0.gds277
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 8.112 48.846 8.312 ;
 END
 END vccd_1p0.gds277
 PIN vccd_1p0.gds278
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 9.0475 49.038 9.2475 ;
 END
 END vccd_1p0.gds278
 PIN vccd_1p0.gds279
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 8.094 49.846 8.294 ;
 END
 END vccd_1p0.gds279
 PIN vccd_1p0.gds280
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 8.094 49.602 8.294 ;
 END
 END vccd_1p0.gds280
 PIN vccd_1p0.gds281
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 8.06 47.002 8.26 ;
 END
 END vccd_1p0.gds281
 PIN vccd_1p0.gds282
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 8.056 46.758 8.256 ;
 END
 END vccd_1p0.gds282
 PIN vccd_1p0.gds283
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 8.0145 46.63 8.2145 ;
 END
 END vccd_1p0.gds283
 PIN vccd_1p0.gds284
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 8.984 50.33 9.184 ;
 END
 END vccd_1p0.gds284
 PIN vccd_1p0.gds285
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 7.724 50.33 7.924 ;
 END
 END vccd_1p0.gds285
 PIN vccd_1p0.gds286
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 6.464 50.33 6.664 ;
 END
 END vccd_1p0.gds286
 PIN vccd_1p0.gds287
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 8.0385 51.678 8.2385 ;
 END
 END vccd_1p0.gds287
 PIN vccd_1p0.gds288
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 8.0145 52.194 8.2145 ;
 END
 END vccd_1p0.gds288
 PIN vccd_1p0.gds289
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 8.056 52.066 8.256 ;
 END
 END vccd_1p0.gds289
 PIN vccd_1p0.gds290
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 7.9635 51.258 8.1635 ;
 END
 END vccd_1p0.gds290
 PIN vccd_1p0.gds291
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 8.06 51.838 8.26 ;
 END
 END vccd_1p0.gds291
 PIN vccd_1p0.gds292
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 8.0185 57.946 8.2185 ;
 END
 END vccd_1p0.gds292
 PIN vccd_1p0.gds293
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 8.92 65.134 9.12 ;
 END
 END vccd_1p0.gds293
 PIN vccd_1p0.gds294
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 10.18 65.134 10.38 ;
 END
 END vccd_1p0.gds294
 PIN vccd_1p0.gds295
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 6.4 65.134 6.6 ;
 END
 END vccd_1p0.gds295
 PIN vccd_1p0.gds296
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 7.66 65.134 7.86 ;
 END
 END vccd_1p0.gds296
 PIN vccd_1p0.gds297
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 7.86 64.894 8.06 ;
 END
 END vccd_1p0.gds297
 PIN vccd_1p0.gds298
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 7.9375 64.294 8.1375 ;
 END
 END vccd_1p0.gds298
 PIN vccd_1p0.gds299
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 8.06 64.054 8.26 ;
 END
 END vccd_1p0.gds299
 PIN vccd_1p0.gds300
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 8.056 63.81 8.256 ;
 END
 END vccd_1p0.gds300
 PIN vccd_1p0.gds301
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 8.0145 63.682 8.2145 ;
 END
 END vccd_1p0.gds301
 PIN vccd_1p0.gds302
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 8.984 67.382 9.184 ;
 END
 END vccd_1p0.gds302
 PIN vccd_1p0.gds303
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 8.92 65.554 9.12 ;
 END
 END vccd_1p0.gds303
 PIN vccd_1p0.gds304
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 7.724 67.382 7.924 ;
 END
 END vccd_1p0.gds304
 PIN vccd_1p0.gds305
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 7.66 65.554 7.86 ;
 END
 END vccd_1p0.gds305
 PIN vccd_1p0.gds306
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 7.7875 66.09 7.9875 ;
 END
 END vccd_1p0.gds306
 PIN vccd_1p0.gds307
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 6.464 67.382 6.664 ;
 END
 END vccd_1p0.gds307
 PIN vccd_1p0.gds308
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 6.4 65.554 6.6 ;
 END
 END vccd_1p0.gds308
 PIN vccd_1p0.gds309
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 6.5275 66.09 6.7275 ;
 END
 END vccd_1p0.gds309
 PIN vccd_1p0.gds310
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 8.112 66.446 8.312 ;
 END
 END vccd_1p0.gds310
 PIN vccd_1p0.gds311
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 10.3005 65.554 10.5005 ;
 END
 END vccd_1p0.gds311
 PIN vccd_1p0.gds312
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 10.4255 66.09 10.6255 ;
 END
 END vccd_1p0.gds312
 PIN vccd_1p0.gds313
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 8.112 65.898 8.312 ;
 END
 END vccd_1p0.gds313
 PIN vccd_1p0.gds314
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 8.0385 68.73 8.2385 ;
 END
 END vccd_1p0.gds314
 PIN vccd_1p0.gds315
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 8.0145 69.246 8.2145 ;
 END
 END vccd_1p0.gds315
 PIN vccd_1p0.gds316
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 9.0475 66.09 9.2475 ;
 END
 END vccd_1p0.gds316
 PIN vccd_1p0.gds317
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 8.056 69.118 8.256 ;
 END
 END vccd_1p0.gds317
 PIN vccd_1p0.gds318
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 7.9635 68.31 8.1635 ;
 END
 END vccd_1p0.gds318
 PIN vccd_1p0.gds319
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 8.094 66.898 8.294 ;
 END
 END vccd_1p0.gds319
 PIN vccd_1p0.gds320
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 8.094 66.654 8.294 ;
 END
 END vccd_1p0.gds320
 PIN vccd_1p0.gds321
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 8.06 68.89 8.26 ;
 END
 END vccd_1p0.gds321
 PIN vccd_1p0.gds322
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 13.669 0.43 13.869 ;
 END
 END vccd_1p0.gds322
 PIN vccd_1p0.gds323
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 13.4415 0.548 13.6415 ;
 END
 END vccd_1p0.gds323
 PIN vccd_1p0.gds324
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 13.1 1.542 13.3 ;
 END
 END vccd_1p0.gds324
 PIN vccd_1p0.gds325
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 13.118 0.858 13.318 ;
 END
 END vccd_1p0.gds325
 PIN vccd_1p0.gds326
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 13.097 1.362 13.297 ;
 END
 END vccd_1p0.gds326
 PIN vccd_1p0.gds327
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 10.923 1.782 11.123 ;
 END
 END vccd_1p0.gds327
 PIN vccd_1p0.gds328
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 13.1235 1.218 13.3235 ;
 END
 END vccd_1p0.gds328
 PIN vccd_1p0.gds329
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 12.9015 1.962 13.1015 ;
 END
 END vccd_1p0.gds329
 PIN vccd_1p0.gds330
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 12.749 2.462 12.949 ;
 END
 END vccd_1p0.gds330
 PIN vccd_1p0.gds331
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 11.037 2.622 11.237 ;
 END
 END vccd_1p0.gds331
 PIN vccd_1p0.gds332
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 13.2055 1.09 13.4055 ;
 END
 END vccd_1p0.gds332
 PIN vccd_1p0.gds333
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 13.117 3.042 13.317 ;
 END
 END vccd_1p0.gds333
 PIN vccd_1p0.gds334
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 13.5 2.882 13.7 ;
 END
 END vccd_1p0.gds334
 PIN vccd_1p0.gds335
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 13.2015 3.262 13.4015 ;
 END
 END vccd_1p0.gds335
 PIN vccd_1p0.gds336
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 11.0805 4.738 11.2805 ;
 END
 END vccd_1p0.gds336
 PIN vccd_1p0.gds337
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 13.1105 3.39 13.3105 ;
 END
 END vccd_1p0.gds337
 PIN vccd_1p0.gds338
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 11.2575 3.666 11.4575 ;
 END
 END vccd_1p0.gds338
 PIN vccd_1p0.gds339
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 11.219 4.066 11.419 ;
 END
 END vccd_1p0.gds339
 PIN vccd_1p0.gds340
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 13.3505 3.858 13.5505 ;
 END
 END vccd_1p0.gds340
 PIN vccd_1p0.gds341
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 13.226 4.546 13.426 ;
 END
 END vccd_1p0.gds341
 PIN vccd_1p0.gds342
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 10.799 4.258 10.999 ;
 END
 END vccd_1p0.gds342
 PIN vccd_1p0.gds343
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 13.469 5.01 13.669 ;
 END
 END vccd_1p0.gds343
 PIN vccd_1p0.gds344
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 12.77 2.622 12.97 ;
 END
 END vccd_1p0.gds344
 PIN vccd_1p0.gds345
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.982 15.158 10.022 15.358 ;
 END
 END vccd_1p0.gds345
 PIN vccd_1p0.gds346
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.31 15.158 9.35 15.358 ;
 END
 END vccd_1p0.gds346
 PIN vccd_1p0.gds347
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.638 15.158 8.678 15.358 ;
 END
 END vccd_1p0.gds347
 PIN vccd_1p0.gds348
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.966 15.158 8.006 15.358 ;
 END
 END vccd_1p0.gds348
 PIN vccd_1p0.gds349
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.294 15.158 7.334 15.358 ;
 END
 END vccd_1p0.gds349
 PIN vccd_1p0.gds350
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.046 11.746 10.086 11.946 ;
 END
 END vccd_1p0.gds350
 PIN vccd_1p0.gds351
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.374 11.746 9.414 11.946 ;
 END
 END vccd_1p0.gds351
 PIN vccd_1p0.gds352
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.702 11.746 8.742 11.946 ;
 END
 END vccd_1p0.gds352
 PIN vccd_1p0.gds353
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.03 11.746 8.07 11.946 ;
 END
 END vccd_1p0.gds353
 PIN vccd_1p0.gds354
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.848 12.7995 9.894 12.9995 ;
 END
 END vccd_1p0.gds354
 PIN vccd_1p0.gds355
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.176 12.7995 9.222 12.9995 ;
 END
 END vccd_1p0.gds355
 PIN vccd_1p0.gds356
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.504 12.7995 8.55 12.9995 ;
 END
 END vccd_1p0.gds356
 PIN vccd_1p0.gds357
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.832 12.7995 7.878 12.9995 ;
 END
 END vccd_1p0.gds357
 PIN vccd_1p0.gds358
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.16 12.821 7.206 13.021 ;
 END
 END vccd_1p0.gds358
 PIN vccd_1p0.gds359
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 12.672 6.838 12.872 ;
 END
 END vccd_1p0.gds359
 PIN vccd_1p0.gds360
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 11.0685 6.05 11.2685 ;
 END
 END vccd_1p0.gds360
 PIN vccd_1p0.gds361
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 10.586 6.306 10.786 ;
 END
 END vccd_1p0.gds361
 PIN vccd_1p0.gds362
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 11.485 5.41 11.685 ;
 END
 END vccd_1p0.gds362
 PIN vccd_1p0.gds363
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 11.167 5.922 11.367 ;
 END
 END vccd_1p0.gds363
 PIN vccd_1p0.gds364
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 13.392 5.602 13.592 ;
 END
 END vccd_1p0.gds364
 PIN vccd_1p0.gds365
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 14.0275 6.306 14.2275 ;
 END
 END vccd_1p0.gds365
 PIN vccd_1p0.gds366
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.358 12.032 7.398 12.232 ;
 END
 END vccd_1p0.gds366
 PIN vccd_1p0.gds367
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 13.2965 6.582 13.4965 ;
 END
 END vccd_1p0.gds367
 PIN vccd_1p0.gds368
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.998 15.158 12.038 15.358 ;
 END
 END vccd_1p0.gds368
 PIN vccd_1p0.gds369
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.326 15.158 11.366 15.358 ;
 END
 END vccd_1p0.gds369
 PIN vccd_1p0.gds370
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.654 15.158 10.694 15.358 ;
 END
 END vccd_1p0.gds370
 PIN vccd_1p0.gds371
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.062 11.7935 12.102 11.9935 ;
 END
 END vccd_1p0.gds371
 PIN vccd_1p0.gds372
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.39 11.746 11.43 11.946 ;
 END
 END vccd_1p0.gds372
 PIN vccd_1p0.gds373
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.718 11.746 10.758 11.946 ;
 END
 END vccd_1p0.gds373
 PIN vccd_1p0.gds374
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 12.6235 14.934 12.8235 ;
 END
 END vccd_1p0.gds374
 PIN vccd_1p0.gds375
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 14.352 13.138 14.552 ;
 END
 END vccd_1p0.gds375
 PIN vccd_1p0.gds376
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 13.2705 15.29 13.4705 ;
 END
 END vccd_1p0.gds376
 PIN vccd_1p0.gds377
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 13.976 12.654 14.176 ;
 END
 END vccd_1p0.gds377
 PIN vccd_1p0.gds378
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.678 12.354 12.718 12.554 ;
 END
 END vccd_1p0.gds378
 PIN vccd_1p0.gds379
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.262 10.933 13.318 11.133 ;
 END
 END vccd_1p0.gds379
 PIN vccd_1p0.gds380
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 11.493 13.978 11.693 ;
 END
 END vccd_1p0.gds380
 PIN vccd_1p0.gds381
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 10.658 13.738 10.858 ;
 END
 END vccd_1p0.gds381
 PIN vccd_1p0.gds382
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 10.8985 14.742 11.0985 ;
 END
 END vccd_1p0.gds382
 PIN vccd_1p0.gds383
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 10.904 12.898 11.104 ;
 END
 END vccd_1p0.gds383
 PIN vccd_1p0.gds384
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 10.657 12.526 10.857 ;
 END
 END vccd_1p0.gds384
 PIN vccd_1p0.gds385
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.864 12.7995 11.91 12.9995 ;
 END
 END vccd_1p0.gds385
 PIN vccd_1p0.gds386
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.192 12.7995 11.238 12.9995 ;
 END
 END vccd_1p0.gds386
 PIN vccd_1p0.gds387
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.52 12.7995 10.566 12.9995 ;
 END
 END vccd_1p0.gds387
 PIN vccd_1p0.gds388
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.894 15.158 19.934 15.358 ;
 END
 END vccd_1p0.gds388
 PIN vccd_1p0.gds389
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.222 15.158 19.262 15.358 ;
 END
 END vccd_1p0.gds389
 PIN vccd_1p0.gds390
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.55 15.158 18.59 15.358 ;
 END
 END vccd_1p0.gds390
 PIN vccd_1p0.gds391
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.958 11.746 19.998 11.946 ;
 END
 END vccd_1p0.gds391
 PIN vccd_1p0.gds392
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.018 12.2845 17.074 12.4845 ;
 END
 END vccd_1p0.gds392
 PIN vccd_1p0.gds393
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.76 12.7995 19.806 12.9995 ;
 END
 END vccd_1p0.gds393
 PIN vccd_1p0.gds394
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 10.648 16.226 10.848 ;
 END
 END vccd_1p0.gds394
 PIN vccd_1p0.gds395
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 10.632 15.29 10.832 ;
 END
 END vccd_1p0.gds395
 PIN vccd_1p0.gds396
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.606 12.687 15.662 12.887 ;
 END
 END vccd_1p0.gds396
 PIN vccd_1p0.gds397
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.25 13.4085 16.31 13.6085 ;
 END
 END vccd_1p0.gds397
 PIN vccd_1p0.gds398
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.438 13.2885 17.494 13.4885 ;
 END
 END vccd_1p0.gds398
 PIN vccd_1p0.gds399
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 10.9105 17.574 11.1105 ;
 END
 END vccd_1p0.gds399
 PIN vccd_1p0.gds400
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 10.8615 15.742 11.0615 ;
 END
 END vccd_1p0.gds400
 PIN vccd_1p0.gds401
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 10.6245 15.498 10.8245 ;
 END
 END vccd_1p0.gds401
 PIN vccd_1p0.gds402
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 11.443 17.734 11.643 ;
 END
 END vccd_1p0.gds402
 PIN vccd_1p0.gds403
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 10.9335 17.154 11.1335 ;
 END
 END vccd_1p0.gds403
 PIN vccd_1p0.gds404
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 14.821 16.57 15.021 ;
 END
 END vccd_1p0.gds404
 PIN vccd_1p0.gds405
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 12.674 18.09 12.874 ;
 END
 END vccd_1p0.gds405
 PIN vccd_1p0.gds406
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 12.882 17.962 13.082 ;
 END
 END vccd_1p0.gds406
 PIN vccd_1p0.gds407
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.416 12.821 18.462 13.021 ;
 END
 END vccd_1p0.gds407
 PIN vccd_1p0.gds408
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.088 12.7995 19.134 12.9995 ;
 END
 END vccd_1p0.gds408
 PIN vccd_1p0.gds409
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.286 11.746 19.326 11.946 ;
 END
 END vccd_1p0.gds409
 PIN vccd_1p0.gds410
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.614 12.032 18.654 12.232 ;
 END
 END vccd_1p0.gds410
 PIN vccd_1p0.gds411
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.018 15.158 25.058 15.358 ;
 END
 END vccd_1p0.gds411
 PIN vccd_1p0.gds412
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.346 15.282 24.386 15.482 ;
 END
 END vccd_1p0.gds412
 PIN vccd_1p0.gds413
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.254 15.158 23.294 15.358 ;
 END
 END vccd_1p0.gds413
 PIN vccd_1p0.gds414
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.582 15.158 22.622 15.358 ;
 END
 END vccd_1p0.gds414
 PIN vccd_1p0.gds415
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.91 15.158 21.95 15.358 ;
 END
 END vccd_1p0.gds415
 PIN vccd_1p0.gds416
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.238 15.158 21.278 15.358 ;
 END
 END vccd_1p0.gds416
 PIN vccd_1p0.gds417
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.566 15.158 20.606 15.358 ;
 END
 END vccd_1p0.gds417
 PIN vccd_1p0.gds418
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.082 11.746 25.122 11.946 ;
 END
 END vccd_1p0.gds418
 PIN vccd_1p0.gds419
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.41 11.7935 24.45 11.9935 ;
 END
 END vccd_1p0.gds419
 PIN vccd_1p0.gds420
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.318 12.032 23.358 12.232 ;
 END
 END vccd_1p0.gds420
 PIN vccd_1p0.gds421
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.646 11.746 22.686 11.946 ;
 END
 END vccd_1p0.gds421
 PIN vccd_1p0.gds422
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.974 11.746 22.014 11.946 ;
 END
 END vccd_1p0.gds422
 PIN vccd_1p0.gds423
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.302 11.746 21.342 11.946 ;
 END
 END vccd_1p0.gds423
 PIN vccd_1p0.gds424
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.63 11.746 20.67 11.946 ;
 END
 END vccd_1p0.gds424
 PIN vccd_1p0.gds425
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.884 12.7995 24.93 12.9995 ;
 END
 END vccd_1p0.gds425
 PIN vccd_1p0.gds426
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.212 12.821 24.258 13.021 ;
 END
 END vccd_1p0.gds426
 PIN vccd_1p0.gds427
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.12 12.888 23.166 13.088 ;
 END
 END vccd_1p0.gds427
 PIN vccd_1p0.gds428
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.448 12.7995 22.494 12.9995 ;
 END
 END vccd_1p0.gds428
 PIN vccd_1p0.gds429
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.776 12.7995 21.822 12.9995 ;
 END
 END vccd_1p0.gds429
 PIN vccd_1p0.gds430
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.104 12.7995 21.15 12.9995 ;
 END
 END vccd_1p0.gds430
 PIN vccd_1p0.gds431
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.432 12.7995 20.478 12.9995 ;
 END
 END vccd_1p0.gds431
 PIN vccd_1p0.gds432
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 12.765 23.842 12.965 ;
 END
 END vccd_1p0.gds432
 PIN vccd_1p0.gds433
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.05 15.158 29.09 15.358 ;
 END
 END vccd_1p0.gds433
 PIN vccd_1p0.gds434
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.378 15.158 28.418 15.358 ;
 END
 END vccd_1p0.gds434
 PIN vccd_1p0.gds435
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.706 15.158 27.746 15.358 ;
 END
 END vccd_1p0.gds435
 PIN vccd_1p0.gds436
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.034 15.158 27.074 15.358 ;
 END
 END vccd_1p0.gds436
 PIN vccd_1p0.gds437
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.362 15.158 26.402 15.358 ;
 END
 END vccd_1p0.gds437
 PIN vccd_1p0.gds438
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.69 15.158 25.73 15.358 ;
 END
 END vccd_1p0.gds438
 PIN vccd_1p0.gds439
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.114 11.7935 29.154 11.9935 ;
 END
 END vccd_1p0.gds439
 PIN vccd_1p0.gds440
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.442 11.746 28.482 11.946 ;
 END
 END vccd_1p0.gds440
 PIN vccd_1p0.gds441
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.77 11.746 27.81 11.946 ;
 END
 END vccd_1p0.gds441
 PIN vccd_1p0.gds442
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.098 11.746 27.138 11.946 ;
 END
 END vccd_1p0.gds442
 PIN vccd_1p0.gds443
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.426 11.746 26.466 11.946 ;
 END
 END vccd_1p0.gds443
 PIN vccd_1p0.gds444
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.754 11.746 25.794 11.946 ;
 END
 END vccd_1p0.gds444
 PIN vccd_1p0.gds445
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.916 12.7995 28.962 12.9995 ;
 END
 END vccd_1p0.gds445
 PIN vccd_1p0.gds446
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.244 12.7995 28.29 12.9995 ;
 END
 END vccd_1p0.gds446
 PIN vccd_1p0.gds447
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.572 12.7995 27.618 12.9995 ;
 END
 END vccd_1p0.gds447
 PIN vccd_1p0.gds448
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.9 12.7995 26.946 12.9995 ;
 END
 END vccd_1p0.gds448
 PIN vccd_1p0.gds449
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.228 12.7995 26.274 12.9995 ;
 END
 END vccd_1p0.gds449
 PIN vccd_1p0.gds450
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.556 12.7995 25.602 12.9995 ;
 END
 END vccd_1p0.gds450
 PIN vccd_1p0.gds451
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 14.352 30.19 14.552 ;
 END
 END vccd_1p0.gds451
 PIN vccd_1p0.gds452
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 13.976 29.706 14.176 ;
 END
 END vccd_1p0.gds452
 PIN vccd_1p0.gds453
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.73 12.354 29.77 12.554 ;
 END
 END vccd_1p0.gds453
 PIN vccd_1p0.gds454
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 10.904 29.95 11.104 ;
 END
 END vccd_1p0.gds454
 PIN vccd_1p0.gds455
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 10.657 29.578 10.857 ;
 END
 END vccd_1p0.gds455
 PIN vccd_1p0.gds456
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 12.6235 31.986 12.8235 ;
 END
 END vccd_1p0.gds456
 PIN vccd_1p0.gds457
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 13.2705 32.342 13.4705 ;
 END
 END vccd_1p0.gds457
 PIN vccd_1p0.gds458
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.49 13.2885 34.546 13.4885 ;
 END
 END vccd_1p0.gds458
 PIN vccd_1p0.gds459
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.314 10.933 30.37 11.133 ;
 END
 END vccd_1p0.gds459
 PIN vccd_1p0.gds460
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 11.493 31.03 11.693 ;
 END
 END vccd_1p0.gds460
 PIN vccd_1p0.gds461
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.658 12.687 32.714 12.887 ;
 END
 END vccd_1p0.gds461
 PIN vccd_1p0.gds462
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 10.648 33.278 10.848 ;
 END
 END vccd_1p0.gds462
 PIN vccd_1p0.gds463
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 10.8615 32.794 11.0615 ;
 END
 END vccd_1p0.gds463
 PIN vccd_1p0.gds464
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 10.632 32.342 10.832 ;
 END
 END vccd_1p0.gds464
 PIN vccd_1p0.gds465
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 10.8985 31.794 11.0985 ;
 END
 END vccd_1p0.gds465
 PIN vccd_1p0.gds466
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 10.952 34.626 11.152 ;
 END
 END vccd_1p0.gds466
 PIN vccd_1p0.gds467
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 12.674 35.142 12.874 ;
 END
 END vccd_1p0.gds467
 PIN vccd_1p0.gds468
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 12.882 35.014 13.082 ;
 END
 END vccd_1p0.gds468
 PIN vccd_1p0.gds469
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 10.658 30.79 10.858 ;
 END
 END vccd_1p0.gds469
 PIN vccd_1p0.gds470
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 10.9335 34.206 11.1335 ;
 END
 END vccd_1p0.gds470
 PIN vccd_1p0.gds471
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.07 12.2845 34.126 12.4845 ;
 END
 END vccd_1p0.gds471
 PIN vccd_1p0.gds472
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 11.3455 34.786 11.5455 ;
 END
 END vccd_1p0.gds472
 PIN vccd_1p0.gds473
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 10.6245 32.55 10.8245 ;
 END
 END vccd_1p0.gds473
 PIN vccd_1p0.gds474
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.302 13.4085 33.362 13.6085 ;
 END
 END vccd_1p0.gds474
 PIN vccd_1p0.gds475
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 14.821 33.622 15.021 ;
 END
 END vccd_1p0.gds475
 PIN vccd_1p0.gds476
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.634 15.158 39.674 15.358 ;
 END
 END vccd_1p0.gds476
 PIN vccd_1p0.gds477
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.962 15.158 39.002 15.358 ;
 END
 END vccd_1p0.gds477
 PIN vccd_1p0.gds478
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.29 15.158 38.33 15.358 ;
 END
 END vccd_1p0.gds478
 PIN vccd_1p0.gds479
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.618 15.158 37.658 15.358 ;
 END
 END vccd_1p0.gds479
 PIN vccd_1p0.gds480
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.946 15.158 36.986 15.358 ;
 END
 END vccd_1p0.gds480
 PIN vccd_1p0.gds481
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.274 15.158 36.314 15.358 ;
 END
 END vccd_1p0.gds481
 PIN vccd_1p0.gds482
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.602 15.158 35.642 15.358 ;
 END
 END vccd_1p0.gds482
 PIN vccd_1p0.gds483
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.698 11.746 39.738 11.946 ;
 END
 END vccd_1p0.gds483
 PIN vccd_1p0.gds484
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.026 11.746 39.066 11.946 ;
 END
 END vccd_1p0.gds484
 PIN vccd_1p0.gds485
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.354 11.746 38.394 11.946 ;
 END
 END vccd_1p0.gds485
 PIN vccd_1p0.gds486
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.682 11.746 37.722 11.946 ;
 END
 END vccd_1p0.gds486
 PIN vccd_1p0.gds487
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.01 11.746 37.05 11.946 ;
 END
 END vccd_1p0.gds487
 PIN vccd_1p0.gds488
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.338 11.746 36.378 11.946 ;
 END
 END vccd_1p0.gds488
 PIN vccd_1p0.gds489
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.468 12.821 35.514 13.021 ;
 END
 END vccd_1p0.gds489
 PIN vccd_1p0.gds490
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.172 12.888 40.218 13.088 ;
 END
 END vccd_1p0.gds490
 PIN vccd_1p0.gds491
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.5 12.7995 39.546 12.9995 ;
 END
 END vccd_1p0.gds491
 PIN vccd_1p0.gds492
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.828 12.7995 38.874 12.9995 ;
 END
 END vccd_1p0.gds492
 PIN vccd_1p0.gds493
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.156 12.7995 38.202 12.9995 ;
 END
 END vccd_1p0.gds493
 PIN vccd_1p0.gds494
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.484 12.7995 37.53 12.9995 ;
 END
 END vccd_1p0.gds494
 PIN vccd_1p0.gds495
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.812 12.7995 36.858 12.9995 ;
 END
 END vccd_1p0.gds495
 PIN vccd_1p0.gds496
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.14 12.7995 36.186 12.9995 ;
 END
 END vccd_1p0.gds496
 PIN vccd_1p0.gds497
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.666 12.032 35.706 12.232 ;
 END
 END vccd_1p0.gds497
 PIN vccd_1p0.gds498
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.758 15.158 44.798 15.358 ;
 END
 END vccd_1p0.gds498
 PIN vccd_1p0.gds499
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.086 15.158 44.126 15.358 ;
 END
 END vccd_1p0.gds499
 PIN vccd_1p0.gds500
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.414 15.158 43.454 15.358 ;
 END
 END vccd_1p0.gds500
 PIN vccd_1p0.gds501
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.742 15.158 42.782 15.358 ;
 END
 END vccd_1p0.gds501
 PIN vccd_1p0.gds502
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.07 15.158 42.11 15.358 ;
 END
 END vccd_1p0.gds502
 PIN vccd_1p0.gds503
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.398 15.282 41.438 15.482 ;
 END
 END vccd_1p0.gds503
 PIN vccd_1p0.gds504
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.306 15.158 40.346 15.358 ;
 END
 END vccd_1p0.gds504
 PIN vccd_1p0.gds505
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.822 11.746 44.862 11.946 ;
 END
 END vccd_1p0.gds505
 PIN vccd_1p0.gds506
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.15 11.746 44.19 11.946 ;
 END
 END vccd_1p0.gds506
 PIN vccd_1p0.gds507
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.478 11.746 43.518 11.946 ;
 END
 END vccd_1p0.gds507
 PIN vccd_1p0.gds508
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.806 11.746 42.846 11.946 ;
 END
 END vccd_1p0.gds508
 PIN vccd_1p0.gds509
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.134 11.746 42.174 11.946 ;
 END
 END vccd_1p0.gds509
 PIN vccd_1p0.gds510
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.462 11.7935 41.502 11.9935 ;
 END
 END vccd_1p0.gds510
 PIN vccd_1p0.gds511
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.37 12.032 40.41 12.232 ;
 END
 END vccd_1p0.gds511
 PIN vccd_1p0.gds512
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.296 12.7995 45.342 12.9995 ;
 END
 END vccd_1p0.gds512
 PIN vccd_1p0.gds513
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.624 12.7995 44.67 12.9995 ;
 END
 END vccd_1p0.gds513
 PIN vccd_1p0.gds514
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.952 12.7995 43.998 12.9995 ;
 END
 END vccd_1p0.gds514
 PIN vccd_1p0.gds515
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.28 12.7995 43.326 12.9995 ;
 END
 END vccd_1p0.gds515
 PIN vccd_1p0.gds516
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.608 12.7995 42.654 12.9995 ;
 END
 END vccd_1p0.gds516
 PIN vccd_1p0.gds517
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.936 12.7995 41.982 12.9995 ;
 END
 END vccd_1p0.gds517
 PIN vccd_1p0.gds518
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.264 12.821 41.31 13.021 ;
 END
 END vccd_1p0.gds518
 PIN vccd_1p0.gds519
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 12.765 40.894 12.965 ;
 END
 END vccd_1p0.gds519
 PIN vccd_1p0.gds520
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.102 15.158 46.142 15.358 ;
 END
 END vccd_1p0.gds520
 PIN vccd_1p0.gds521
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.43 15.158 45.47 15.358 ;
 END
 END vccd_1p0.gds521
 PIN vccd_1p0.gds522
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 12.6235 49.038 12.8235 ;
 END
 END vccd_1p0.gds522
 PIN vccd_1p0.gds523
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 14.352 47.242 14.552 ;
 END
 END vccd_1p0.gds523
 PIN vccd_1p0.gds524
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 13.2705 49.394 13.4705 ;
 END
 END vccd_1p0.gds524
 PIN vccd_1p0.gds525
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 13.976 46.758 14.176 ;
 END
 END vccd_1p0.gds525
 PIN vccd_1p0.gds526
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.166 11.7935 46.206 11.9935 ;
 END
 END vccd_1p0.gds526
 PIN vccd_1p0.gds527
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.494 11.746 45.534 11.946 ;
 END
 END vccd_1p0.gds527
 PIN vccd_1p0.gds528
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.968 12.7995 46.014 12.9995 ;
 END
 END vccd_1p0.gds528
 PIN vccd_1p0.gds529
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.782 12.354 46.822 12.554 ;
 END
 END vccd_1p0.gds529
 PIN vccd_1p0.gds530
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 10.658 47.842 10.858 ;
 END
 END vccd_1p0.gds530
 PIN vccd_1p0.gds531
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.366 10.933 47.422 11.133 ;
 END
 END vccd_1p0.gds531
 PIN vccd_1p0.gds532
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 11.493 48.082 11.693 ;
 END
 END vccd_1p0.gds532
 PIN vccd_1p0.gds533
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.71 12.687 49.766 12.887 ;
 END
 END vccd_1p0.gds533
 PIN vccd_1p0.gds534
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 10.632 49.394 10.832 ;
 END
 END vccd_1p0.gds534
 PIN vccd_1p0.gds535
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 10.8985 48.846 11.0985 ;
 END
 END vccd_1p0.gds535
 PIN vccd_1p0.gds536
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 10.8615 49.846 11.0615 ;
 END
 END vccd_1p0.gds536
 PIN vccd_1p0.gds537
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 10.6245 49.602 10.8245 ;
 END
 END vccd_1p0.gds537
 PIN vccd_1p0.gds538
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 10.904 47.002 11.104 ;
 END
 END vccd_1p0.gds538
 PIN vccd_1p0.gds539
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 10.657 46.63 10.857 ;
 END
 END vccd_1p0.gds539
 PIN vccd_1p0.gds540
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.67 15.158 54.71 15.358 ;
 END
 END vccd_1p0.gds540
 PIN vccd_1p0.gds541
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.998 15.158 54.038 15.358 ;
 END
 END vccd_1p0.gds541
 PIN vccd_1p0.gds542
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.326 15.158 53.366 15.358 ;
 END
 END vccd_1p0.gds542
 PIN vccd_1p0.gds543
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.654 15.158 52.694 15.358 ;
 END
 END vccd_1p0.gds543
 PIN vccd_1p0.gds544
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.354 13.4085 50.414 13.6085 ;
 END
 END vccd_1p0.gds544
 PIN vccd_1p0.gds545
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.542 13.2885 51.598 13.4885 ;
 END
 END vccd_1p0.gds545
 PIN vccd_1p0.gds546
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 14.821 50.674 15.021 ;
 END
 END vccd_1p0.gds546
 PIN vccd_1p0.gds547
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.52 12.821 52.566 13.021 ;
 END
 END vccd_1p0.gds547
 PIN vccd_1p0.gds548
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.208 12.7995 55.254 12.9995 ;
 END
 END vccd_1p0.gds548
 PIN vccd_1p0.gds549
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.536 12.7995 54.582 12.9995 ;
 END
 END vccd_1p0.gds549
 PIN vccd_1p0.gds550
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.734 11.746 54.774 11.946 ;
 END
 END vccd_1p0.gds550
 PIN vccd_1p0.gds551
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.864 12.7995 53.91 12.9995 ;
 END
 END vccd_1p0.gds551
 PIN vccd_1p0.gds552
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.062 11.746 54.102 11.946 ;
 END
 END vccd_1p0.gds552
 PIN vccd_1p0.gds553
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 10.648 50.33 10.848 ;
 END
 END vccd_1p0.gds553
 PIN vccd_1p0.gds554
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 10.9105 51.678 11.1105 ;
 END
 END vccd_1p0.gds554
 PIN vccd_1p0.gds555
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 12.674 52.194 12.874 ;
 END
 END vccd_1p0.gds555
 PIN vccd_1p0.gds556
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 12.882 52.066 13.082 ;
 END
 END vccd_1p0.gds556
 PIN vccd_1p0.gds557
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 10.9335 51.258 11.1335 ;
 END
 END vccd_1p0.gds557
 PIN vccd_1p0.gds558
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 11.443 51.838 11.643 ;
 END
 END vccd_1p0.gds558
 PIN vccd_1p0.gds559
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.122 12.2845 51.178 12.4845 ;
 END
 END vccd_1p0.gds559
 PIN vccd_1p0.gds560
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.192 12.7995 53.238 12.9995 ;
 END
 END vccd_1p0.gds560
 PIN vccd_1p0.gds561
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.39 11.746 53.43 11.946 ;
 END
 END vccd_1p0.gds561
 PIN vccd_1p0.gds562
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.718 12.032 52.758 12.232 ;
 END
 END vccd_1p0.gds562
 PIN vccd_1p0.gds563
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.358 15.158 57.398 15.358 ;
 END
 END vccd_1p0.gds563
 PIN vccd_1p0.gds564
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.794 15.158 59.834 15.358 ;
 END
 END vccd_1p0.gds564
 PIN vccd_1p0.gds565
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.122 15.158 59.162 15.358 ;
 END
 END vccd_1p0.gds565
 PIN vccd_1p0.gds566
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.45 15.282 58.49 15.482 ;
 END
 END vccd_1p0.gds566
 PIN vccd_1p0.gds567
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.686 15.158 56.726 15.358 ;
 END
 END vccd_1p0.gds567
 PIN vccd_1p0.gds568
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.014 15.158 56.054 15.358 ;
 END
 END vccd_1p0.gds568
 PIN vccd_1p0.gds569
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.342 15.158 55.382 15.358 ;
 END
 END vccd_1p0.gds569
 PIN vccd_1p0.gds570
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.66 12.7995 59.706 12.9995 ;
 END
 END vccd_1p0.gds570
 PIN vccd_1p0.gds571
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.858 11.746 59.898 11.946 ;
 END
 END vccd_1p0.gds571
 PIN vccd_1p0.gds572
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.988 12.7995 59.034 12.9995 ;
 END
 END vccd_1p0.gds572
 PIN vccd_1p0.gds573
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.186 11.746 59.226 11.946 ;
 END
 END vccd_1p0.gds573
 PIN vccd_1p0.gds574
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.316 12.821 58.362 13.021 ;
 END
 END vccd_1p0.gds574
 PIN vccd_1p0.gds575
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.514 11.7935 58.554 11.9935 ;
 END
 END vccd_1p0.gds575
 PIN vccd_1p0.gds576
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.224 12.888 57.27 13.088 ;
 END
 END vccd_1p0.gds576
 PIN vccd_1p0.gds577
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.422 12.032 57.462 12.232 ;
 END
 END vccd_1p0.gds577
 PIN vccd_1p0.gds578
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.552 12.7995 56.598 12.9995 ;
 END
 END vccd_1p0.gds578
 PIN vccd_1p0.gds579
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.75 11.746 56.79 11.946 ;
 END
 END vccd_1p0.gds579
 PIN vccd_1p0.gds580
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.88 12.7995 55.926 12.9995 ;
 END
 END vccd_1p0.gds580
 PIN vccd_1p0.gds581
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.078 11.746 56.118 11.946 ;
 END
 END vccd_1p0.gds581
 PIN vccd_1p0.gds582
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.406 11.746 55.446 11.946 ;
 END
 END vccd_1p0.gds582
 PIN vccd_1p0.gds583
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 12.765 57.946 12.965 ;
 END
 END vccd_1p0.gds583
 PIN vccd_1p0.gds584
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.154 15.158 63.194 15.358 ;
 END
 END vccd_1p0.gds584
 PIN vccd_1p0.gds585
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.482 15.158 62.522 15.358 ;
 END
 END vccd_1p0.gds585
 PIN vccd_1p0.gds586
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.81 15.158 61.85 15.358 ;
 END
 END vccd_1p0.gds586
 PIN vccd_1p0.gds587
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.138 15.158 61.178 15.358 ;
 END
 END vccd_1p0.gds587
 PIN vccd_1p0.gds588
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.466 15.158 60.506 15.358 ;
 END
 END vccd_1p0.gds588
 PIN vccd_1p0.gds589
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 14.352 64.294 14.552 ;
 END
 END vccd_1p0.gds589
 PIN vccd_1p0.gds590
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 13.976 63.81 14.176 ;
 END
 END vccd_1p0.gds590
 PIN vccd_1p0.gds591
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.834 12.354 63.874 12.554 ;
 END
 END vccd_1p0.gds591
 PIN vccd_1p0.gds592
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.02 12.7995 63.066 12.9995 ;
 END
 END vccd_1p0.gds592
 PIN vccd_1p0.gds593
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.218 11.7935 63.258 11.9935 ;
 END
 END vccd_1p0.gds593
 PIN vccd_1p0.gds594
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.348 12.7995 62.394 12.9995 ;
 END
 END vccd_1p0.gds594
 PIN vccd_1p0.gds595
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.546 11.746 62.586 11.946 ;
 END
 END vccd_1p0.gds595
 PIN vccd_1p0.gds596
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.676 12.7995 61.722 12.9995 ;
 END
 END vccd_1p0.gds596
 PIN vccd_1p0.gds597
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.874 11.746 61.914 11.946 ;
 END
 END vccd_1p0.gds597
 PIN vccd_1p0.gds598
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.004 12.7995 61.05 12.9995 ;
 END
 END vccd_1p0.gds598
 PIN vccd_1p0.gds599
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.202 11.746 61.242 11.946 ;
 END
 END vccd_1p0.gds599
 PIN vccd_1p0.gds600
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.332 12.7995 60.378 12.9995 ;
 END
 END vccd_1p0.gds600
 PIN vccd_1p0.gds601
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.53 11.746 60.57 11.946 ;
 END
 END vccd_1p0.gds601
 PIN vccd_1p0.gds602
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 10.658 64.894 10.858 ;
 END
 END vccd_1p0.gds602
 PIN vccd_1p0.gds603
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.418 10.933 64.474 11.133 ;
 END
 END vccd_1p0.gds603
 PIN vccd_1p0.gds604
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 11.493 65.134 11.693 ;
 END
 END vccd_1p0.gds604
 PIN vccd_1p0.gds605
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 10.904 64.054 11.104 ;
 END
 END vccd_1p0.gds605
 PIN vccd_1p0.gds606
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 10.657 63.682 10.857 ;
 END
 END vccd_1p0.gds606
 PIN vccd_1p0.gds607
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.706 15.158 69.746 15.358 ;
 END
 END vccd_1p0.gds607
 PIN vccd_1p0.gds608
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 12.6235 66.09 12.8235 ;
 END
 END vccd_1p0.gds608
 PIN vccd_1p0.gds609
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 13.2705 66.446 13.4705 ;
 END
 END vccd_1p0.gds609
 PIN vccd_1p0.gds610
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.762 12.687 66.818 12.887 ;
 END
 END vccd_1p0.gds610
 PIN vccd_1p0.gds611
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.406 13.4085 67.466 13.6085 ;
 END
 END vccd_1p0.gds611
 PIN vccd_1p0.gds612
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.572 12.821 69.618 13.021 ;
 END
 END vccd_1p0.gds612
 PIN vccd_1p0.gds613
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 10.648 67.382 10.848 ;
 END
 END vccd_1p0.gds613
 PIN vccd_1p0.gds614
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 10.632 66.446 10.832 ;
 END
 END vccd_1p0.gds614
 PIN vccd_1p0.gds615
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 10.8985 65.898 11.0985 ;
 END
 END vccd_1p0.gds615
 PIN vccd_1p0.gds616
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 10.9105 68.73 11.1105 ;
 END
 END vccd_1p0.gds616
 PIN vccd_1p0.gds617
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 12.674 69.246 12.874 ;
 END
 END vccd_1p0.gds617
 PIN vccd_1p0.gds618
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 12.882 69.118 13.082 ;
 END
 END vccd_1p0.gds618
 PIN vccd_1p0.gds619
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 10.9335 68.31 11.1335 ;
 END
 END vccd_1p0.gds619
 PIN vccd_1p0.gds620
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 10.8615 66.898 11.0615 ;
 END
 END vccd_1p0.gds620
 PIN vccd_1p0.gds621
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 10.6245 66.654 10.8245 ;
 END
 END vccd_1p0.gds621
 PIN vccd_1p0.gds622
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 11.443 68.89 11.643 ;
 END
 END vccd_1p0.gds622
 PIN vccd_1p0.gds623
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.174 12.2845 68.23 12.4845 ;
 END
 END vccd_1p0.gds623
 PIN vccd_1p0.gds624
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.244 12.7995 70.29 12.9995 ;
 END
 END vccd_1p0.gds624
 PIN vccd_1p0.gds625
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.77 12.032 69.81 12.232 ;
 END
 END vccd_1p0.gds625
 PIN vccd_1p0.gds626
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.594 13.2885 68.65 13.4885 ;
 END
 END vccd_1p0.gds626
 PIN vccd_1p0.gds627
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 14.821 67.726 15.021 ;
 END
 END vccd_1p0.gds627
 PIN vccd_1p0.gds628
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.41 15.158 74.45 15.358 ;
 END
 END vccd_1p0.gds628
 PIN vccd_1p0.gds629
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.738 15.158 73.778 15.358 ;
 END
 END vccd_1p0.gds629
 PIN vccd_1p0.gds630
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.066 15.158 73.106 15.358 ;
 END
 END vccd_1p0.gds630
 PIN vccd_1p0.gds631
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.394 15.158 72.434 15.358 ;
 END
 END vccd_1p0.gds631
 PIN vccd_1p0.gds632
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.722 15.158 71.762 15.358 ;
 END
 END vccd_1p0.gds632
 PIN vccd_1p0.gds633
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.05 15.158 71.09 15.358 ;
 END
 END vccd_1p0.gds633
 PIN vccd_1p0.gds634
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.378 15.158 70.418 15.358 ;
 END
 END vccd_1p0.gds634
 PIN vccd_1p0.gds635
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.276 12.924 74.322 13.124 ;
 END
 END vccd_1p0.gds635
 PIN vccd_1p0.gds636
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.474 11.746 74.514 11.946 ;
 END
 END vccd_1p0.gds636
 PIN vccd_1p0.gds637
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.604 12.7995 73.65 12.9995 ;
 END
 END vccd_1p0.gds637
 PIN vccd_1p0.gds638
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.802 11.746 73.842 11.946 ;
 END
 END vccd_1p0.gds638
 PIN vccd_1p0.gds639
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.932 12.7995 72.978 12.9995 ;
 END
 END vccd_1p0.gds639
 PIN vccd_1p0.gds640
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.13 11.746 73.17 11.946 ;
 END
 END vccd_1p0.gds640
 PIN vccd_1p0.gds641
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.26 12.7995 72.306 12.9995 ;
 END
 END vccd_1p0.gds641
 PIN vccd_1p0.gds642
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.458 11.746 72.498 11.946 ;
 END
 END vccd_1p0.gds642
 PIN vccd_1p0.gds643
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.588 12.7995 71.634 12.9995 ;
 END
 END vccd_1p0.gds643
 PIN vccd_1p0.gds644
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.786 11.746 71.826 11.946 ;
 END
 END vccd_1p0.gds644
 PIN vccd_1p0.gds645
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.916 12.7995 70.962 12.9995 ;
 END
 END vccd_1p0.gds645
 PIN vccd_1p0.gds646
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.114 11.746 71.154 11.946 ;
 END
 END vccd_1p0.gds646
 PIN vccd_1p0.gds647
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.442 11.746 70.482 11.946 ;
 END
 END vccd_1p0.gds647
 PIN vccd_1p0.gds648
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 19.0995 0.43 19.2995 ;
 END
 END vccd_1p0.gds648
 PIN vccd_1p0.gds649
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 19.157 1.542 19.357 ;
 END
 END vccd_1p0.gds649
 PIN vccd_1p0.gds650
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 17.897 0.548 18.097 ;
 END
 END vccd_1p0.gds650
 PIN vccd_1p0.gds651
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 17.1195 1.542 17.3195 ;
 END
 END vccd_1p0.gds651
 PIN vccd_1p0.gds652
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 20.417 1.542 20.617 ;
 END
 END vccd_1p0.gds652
 PIN vccd_1p0.gds653
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 20.2995 5.202 20.4995 ;
 END
 END vccd_1p0.gds653
 PIN vccd_1p0.gds654
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 18.126 0.858 18.326 ;
 END
 END vccd_1p0.gds654
 PIN vccd_1p0.gds655
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 17.803 1.362 18.003 ;
 END
 END vccd_1p0.gds655
 PIN vccd_1p0.gds656
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 17.8815 1.218 18.0815 ;
 END
 END vccd_1p0.gds656
 PIN vccd_1p0.gds657
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 18.0525 1.09 18.2525 ;
 END
 END vccd_1p0.gds657
 PIN vccd_1p0.gds658
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 16.632 2.462 16.832 ;
 END
 END vccd_1p0.gds658
 PIN vccd_1p0.gds659
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 19.341 1.782 19.541 ;
 END
 END vccd_1p0.gds659
 PIN vccd_1p0.gds660
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 19.848 2.202 20.048 ;
 END
 END vccd_1p0.gds660
 PIN vccd_1p0.gds661
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 17.573 2.622 17.773 ;
 END
 END vccd_1p0.gds661
 PIN vccd_1p0.gds662
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 20.3165 2.462 20.5165 ;
 END
 END vccd_1p0.gds662
 PIN vccd_1p0.gds663
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 17.4035 1.962 17.6035 ;
 END
 END vccd_1p0.gds663
 PIN vccd_1p0.gds664
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 17.787 3.042 17.987 ;
 END
 END vccd_1p0.gds664
 PIN vccd_1p0.gds665
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 18.532 5.202 18.732 ;
 END
 END vccd_1p0.gds665
 PIN vccd_1p0.gds666
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 17.8705 2.882 18.0705 ;
 END
 END vccd_1p0.gds666
 PIN vccd_1p0.gds667
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 18.039 3.262 18.239 ;
 END
 END vccd_1p0.gds667
 PIN vccd_1p0.gds668
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 17.763 3.39 17.963 ;
 END
 END vccd_1p0.gds668
 PIN vccd_1p0.gds669
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 17.925 3.858 18.125 ;
 END
 END vccd_1p0.gds669
 PIN vccd_1p0.gds670
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 16.732 4.258 16.932 ;
 END
 END vccd_1p0.gds670
 PIN vccd_1p0.gds671
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 17.737 4.546 17.937 ;
 END
 END vccd_1p0.gds671
 PIN vccd_1p0.gds672
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 17.696 5.01 17.896 ;
 END
 END vccd_1p0.gds672
 PIN vccd_1p0.gds673
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 3.584 19.1835 3.64 19.3835 ;
 RECT 3.584 20.4435 3.64 20.6435 ;
 RECT 4.34 19.282 4.396 19.482 ;
 RECT 4.172 19.282 4.228 19.482 ;
 RECT 4.76 19.2415 4.816 19.4415 ;
 RECT 5.096 19.282 5.152 19.482 ;
 RECT 4.928 19.2415 4.984 19.4415 ;
 END
 END vccd_1p0.gds673
 PIN vccd_1p0.gds674
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.566 15.7365 9.606 15.9365 ;
 END
 END vccd_1p0.gds674
 PIN vccd_1p0.gds675
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.894 15.7365 8.934 15.9365 ;
 END
 END vccd_1p0.gds675
 PIN vccd_1p0.gds676
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.222 15.7365 8.262 15.9365 ;
 END
 END vccd_1p0.gds676
 PIN vccd_1p0.gds677
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.55 15.7365 7.59 15.9365 ;
 END
 END vccd_1p0.gds677
 PIN vccd_1p0.gds678
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.798 17.5755 9.858 17.7755 ;
 END
 END vccd_1p0.gds678
 PIN vccd_1p0.gds679
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.134 17.544 10.194 17.744 ;
 END
 END vccd_1p0.gds679
 PIN vccd_1p0.gds680
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.126 17.5755 9.186 17.7755 ;
 END
 END vccd_1p0.gds680
 PIN vccd_1p0.gds681
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.462 17.544 9.522 17.744 ;
 END
 END vccd_1p0.gds681
 PIN vccd_1p0.gds682
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.454 17.5755 8.514 17.7755 ;
 END
 END vccd_1p0.gds682
 PIN vccd_1p0.gds683
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.79 17.544 8.85 17.744 ;
 END
 END vccd_1p0.gds683
 PIN vccd_1p0.gds684
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.782 17.5755 7.842 17.7755 ;
 END
 END vccd_1p0.gds684
 PIN vccd_1p0.gds685
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.118 17.544 8.178 17.744 ;
 END
 END vccd_1p0.gds685
 PIN vccd_1p0.gds686
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.11 17.5755 7.17 17.7755 ;
 END
 END vccd_1p0.gds686
 PIN vccd_1p0.gds687
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.446 17.544 7.506 17.744 ;
 END
 END vccd_1p0.gds687
 PIN vccd_1p0.gds688
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 17.9975 6.838 18.1975 ;
 END
 END vccd_1p0.gds688
 PIN vccd_1p0.gds689
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 20.323 6.05 20.523 ;
 END
 END vccd_1p0.gds689
 PIN vccd_1p0.gds690
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 16.007 5.41 16.207 ;
 END
 END vccd_1p0.gds690
 PIN vccd_1p0.gds691
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 19.5705 5.922 19.7705 ;
 END
 END vccd_1p0.gds691
 PIN vccd_1p0.gds692
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 17.8405 5.602 18.0405 ;
 END
 END vccd_1p0.gds692
 PIN vccd_1p0.gds693
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 18.7425 6.306 18.9425 ;
 END
 END vccd_1p0.gds693
 PIN vccd_1p0.gds694
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 17.9025 6.582 18.1025 ;
 END
 END vccd_1p0.gds694
 PIN vccd_1p0.gds695
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 9.968 18.0955 10.024 18.2955 ;
 RECT 9.8 18.0655 9.856 18.2655 ;
 RECT 9.296 18.0955 9.352 18.2955 ;
 RECT 9.128 18.0655 9.184 18.2655 ;
 RECT 9.632 17.964 9.688 18.164 ;
 RECT 8.624 18.0955 8.68 18.2955 ;
 RECT 8.456 18.0655 8.512 18.2655 ;
 RECT 8.96 17.964 9.016 18.164 ;
 RECT 7.952 18.0955 8.008 18.2955 ;
 RECT 7.784 18.0655 7.84 18.2655 ;
 RECT 8.288 17.964 8.344 18.164 ;
 RECT 6.944 17.964 7 18.164 ;
 RECT 7.28 18.0955 7.336 18.2955 ;
 RECT 7.112 18.0655 7.168 18.2655 ;
 RECT 7.616 17.964 7.672 18.164 ;
 RECT 5.6 19.282 5.656 19.482 ;
 RECT 5.432 19.1935 5.488 19.3935 ;
 RECT 5.264 19.282 5.32 19.482 ;
 RECT 5.936 19.1935 5.992 19.3935 ;
 RECT 5.768 19.1935 5.824 19.3935 ;
 RECT 6.44 19.2105 6.496 19.4105 ;
 RECT 6.272 19.1935 6.328 19.3935 ;
 RECT 6.104 19.282 6.16 19.482 ;
 END
 END vccd_1p0.gds695
 PIN vccd_1p0.gds696
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 19.504 13.978 19.704 ;
 END
 END vccd_1p0.gds696
 PIN vccd_1p0.gds697
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.582 15.7365 11.622 15.9365 ;
 END
 END vccd_1p0.gds697
 PIN vccd_1p0.gds698
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.91 15.7365 10.95 15.9365 ;
 END
 END vccd_1p0.gds698
 PIN vccd_1p0.gds699
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.238 15.7365 10.278 15.9365 ;
 END
 END vccd_1p0.gds699
 PIN vccd_1p0.gds700
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 17.697 14.398 17.897 ;
 END
 END vccd_1p0.gds700
 PIN vccd_1p0.gds701
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 19.504 14.398 19.704 ;
 END
 END vccd_1p0.gds701
 PIN vccd_1p0.gds702
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 18.5525 13.738 18.7525 ;
 END
 END vccd_1p0.gds702
 PIN vccd_1p0.gds703
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 18.995 13.138 19.195 ;
 END
 END vccd_1p0.gds703
 PIN vccd_1p0.gds704
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 17.3415 12.898 17.5415 ;
 END
 END vccd_1p0.gds704
 PIN vccd_1p0.gds705
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 18.271 13.978 18.471 ;
 END
 END vccd_1p0.gds705
 PIN vccd_1p0.gds706
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 15.453 13.978 15.653 ;
 END
 END vccd_1p0.gds706
 PIN vccd_1p0.gds707
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 16.607 14.934 16.807 ;
 END
 END vccd_1p0.gds707
 PIN vccd_1p0.gds708
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.254 15.7405 12.294 15.9405 ;
 END
 END vccd_1p0.gds708
 PIN vccd_1p0.gds709
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 16.7735 14.742 16.9735 ;
 END
 END vccd_1p0.gds709
 PIN vccd_1p0.gds710
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 19.6315 14.934 19.8315 ;
 END
 END vccd_1p0.gds710
 PIN vccd_1p0.gds711
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.814 17.5755 11.874 17.7755 ;
 END
 END vccd_1p0.gds711
 PIN vccd_1p0.gds712
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.15 17.544 12.21 17.744 ;
 END
 END vccd_1p0.gds712
 PIN vccd_1p0.gds713
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.142 17.5755 11.202 17.7755 ;
 END
 END vccd_1p0.gds713
 PIN vccd_1p0.gds714
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.478 17.544 11.538 17.744 ;
 END
 END vccd_1p0.gds714
 PIN vccd_1p0.gds715
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.47 17.5755 10.53 17.7755 ;
 END
 END vccd_1p0.gds715
 PIN vccd_1p0.gds716
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.806 17.544 10.866 17.744 ;
 END
 END vccd_1p0.gds716
 PIN vccd_1p0.gds717
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 18.0675 12.654 18.2675 ;
 END
 END vccd_1p0.gds717
 PIN vccd_1p0.gds718
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 12.992 16.967 13.048 17.167 ;
 RECT 12.74 17.5945 12.796 17.7945 ;
 RECT 13.244 17.47 13.3 17.67 ;
 RECT 12.572 17.666 12.628 17.866 ;
 RECT 15.092 17.774 15.148 17.974 ;
 RECT 14.924 17.774 14.98 17.974 ;
 RECT 14.756 17.666 14.812 17.866 ;
 RECT 14.588 17.5945 14.644 17.7945 ;
 RECT 14.42 17.5945 14.476 17.7945 ;
 RECT 14.252 17.5945 14.308 17.7945 ;
 RECT 14.084 17.774 14.14 17.974 ;
 RECT 13.916 17.774 13.972 17.974 ;
 RECT 13.748 17.666 13.804 17.866 ;
 RECT 11.984 18.0955 12.04 18.2955 ;
 RECT 11.816 18.0655 11.872 18.2655 ;
 RECT 12.32 17.964 12.376 18.164 ;
 RECT 11.312 18.0955 11.368 18.2955 ;
 RECT 11.144 18.0655 11.2 18.2655 ;
 RECT 11.648 17.964 11.704 18.164 ;
 RECT 10.64 18.0955 10.696 18.2955 ;
 RECT 10.472 18.0655 10.528 18.2655 ;
 RECT 10.976 17.964 11.032 18.164 ;
 RECT 10.304 17.964 10.36 18.164 ;
 END
 END vccd_1p0.gds718
 PIN vccd_1p0.gds719
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.15 15.7365 20.19 15.9365 ;
 END
 END vccd_1p0.gds719
 PIN vccd_1p0.gds720
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.478 15.7365 19.518 15.9365 ;
 END
 END vccd_1p0.gds720
 PIN vccd_1p0.gds721
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.71 17.5755 19.77 17.7755 ;
 END
 END vccd_1p0.gds721
 PIN vccd_1p0.gds722
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.046 17.544 20.106 17.744 ;
 END
 END vccd_1p0.gds722
 PIN vccd_1p0.gds723
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.334 17.795 16.39 17.995 ;
 END
 END vccd_1p0.gds723
 PIN vccd_1p0.gds724
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 19.568 16.226 19.768 ;
 END
 END vccd_1p0.gds724
 PIN vccd_1p0.gds725
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 18.2 15.742 18.4 ;
 END
 END vccd_1p0.gds725
 PIN vccd_1p0.gds726
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 17.1315 16.226 17.3315 ;
 END
 END vccd_1p0.gds726
 PIN vccd_1p0.gds727
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 19.436 15.29 19.636 ;
 END
 END vccd_1p0.gds727
 PIN vccd_1p0.gds728
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 15.8895 18.09 16.0895 ;
 END
 END vccd_1p0.gds728
 PIN vccd_1p0.gds729
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 15.902 17.962 16.102 ;
 END
 END vccd_1p0.gds729
 PIN vccd_1p0.gds730
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 19.599 18.09 19.799 ;
 END
 END vccd_1p0.gds730
 PIN vccd_1p0.gds731
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 19.4835 17.962 19.6835 ;
 END
 END vccd_1p0.gds731
 PIN vccd_1p0.gds732
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 17.9255 15.498 18.1255 ;
 END
 END vccd_1p0.gds732
 PIN vccd_1p0.gds733
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 19.3655 17.734 19.5655 ;
 END
 END vccd_1p0.gds733
 PIN vccd_1p0.gds734
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 17.4875 17.574 17.6875 ;
 END
 END vccd_1p0.gds734
 PIN vccd_1p0.gds735
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 17.143 17.154 17.343 ;
 END
 END vccd_1p0.gds735
 PIN vccd_1p0.gds736
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.038 17.5755 19.098 17.7755 ;
 END
 END vccd_1p0.gds736
 PIN vccd_1p0.gds737
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.374 17.544 19.434 17.744 ;
 END
 END vccd_1p0.gds737
 PIN vccd_1p0.gds738
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.366 17.4515 18.426 17.6515 ;
 END
 END vccd_1p0.gds738
 PIN vccd_1p0.gds739
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.702 17.544 18.762 17.744 ;
 END
 END vccd_1p0.gds739
 PIN vccd_1p0.gds740
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.806 15.7365 18.846 15.9365 ;
 END
 END vccd_1p0.gds740
 PIN vccd_1p0.gds741
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 19.88 18.0955 19.936 18.2955 ;
 RECT 19.712 18.0655 19.768 18.2655 ;
 RECT 20.216 17.964 20.272 18.164 ;
 RECT 15.26 17.68 15.316 17.88 ;
 RECT 16.772 17.4835 16.828 17.6835 ;
 RECT 16.604 17.4835 16.66 17.6835 ;
 RECT 16.436 17.4835 16.492 17.6835 ;
 RECT 16.268 17.4835 16.324 17.6835 ;
 RECT 16.1 17.4835 16.156 17.6835 ;
 RECT 15.932 17.4835 15.988 17.6835 ;
 RECT 15.764 17.4835 15.82 17.6835 ;
 RECT 15.428 17.68 15.484 17.88 ;
 RECT 16.94 17.4835 16.996 17.6835 ;
 RECT 17.276 17.68 17.332 17.88 ;
 RECT 17.108 17.68 17.164 17.88 ;
 RECT 15.596 17.5945 15.652 17.7945 ;
 RECT 17.612 17.5945 17.668 17.7945 ;
 RECT 17.444 17.5945 17.5 17.7945 ;
 RECT 17.948 17.4975 18.004 17.6975 ;
 RECT 19.208 18.0955 19.264 18.2955 ;
 RECT 19.04 18.0655 19.096 18.2655 ;
 RECT 19.544 17.964 19.6 18.164 ;
 RECT 18.536 18.0955 18.592 18.2955 ;
 RECT 18.2 17.964 18.256 18.164 ;
 RECT 18.368 18.0655 18.424 18.2655 ;
 RECT 18.872 17.964 18.928 18.164 ;
 RECT 17.78 17.68 17.836 17.88 ;
 END
 END vccd_1p0.gds741
 PIN vccd_1p0.gds742
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.838 15.7365 22.878 15.9365 ;
 END
 END vccd_1p0.gds742
 PIN vccd_1p0.gds743
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.166 15.7365 22.206 15.9365 ;
 END
 END vccd_1p0.gds743
 PIN vccd_1p0.gds744
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.494 15.7365 21.534 15.9365 ;
 END
 END vccd_1p0.gds744
 PIN vccd_1p0.gds745
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.822 15.7365 20.862 15.9365 ;
 END
 END vccd_1p0.gds745
 PIN vccd_1p0.gds746
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.834 17.5755 24.894 17.7755 ;
 END
 END vccd_1p0.gds746
 PIN vccd_1p0.gds747
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.17 17.544 25.23 17.744 ;
 END
 END vccd_1p0.gds747
 PIN vccd_1p0.gds748
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.162 17.5755 24.222 17.7755 ;
 END
 END vccd_1p0.gds748
 PIN vccd_1p0.gds749
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.498 17.544 24.558 17.744 ;
 END
 END vccd_1p0.gds749
 PIN vccd_1p0.gds750
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.07 17.5755 23.13 17.7755 ;
 END
 END vccd_1p0.gds750
 PIN vccd_1p0.gds751
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.406 17.544 23.466 17.744 ;
 END
 END vccd_1p0.gds751
 PIN vccd_1p0.gds752
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.398 17.5755 22.458 17.7755 ;
 END
 END vccd_1p0.gds752
 PIN vccd_1p0.gds753
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.734 17.544 22.794 17.744 ;
 END
 END vccd_1p0.gds753
 PIN vccd_1p0.gds754
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.726 17.5755 21.786 17.7755 ;
 END
 END vccd_1p0.gds754
 PIN vccd_1p0.gds755
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.062 17.544 22.122 17.744 ;
 END
 END vccd_1p0.gds755
 PIN vccd_1p0.gds756
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.054 17.5755 21.114 17.7755 ;
 END
 END vccd_1p0.gds756
 PIN vccd_1p0.gds757
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.39 17.544 21.45 17.744 ;
 END
 END vccd_1p0.gds757
 PIN vccd_1p0.gds758
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.382 17.5755 20.442 17.7755 ;
 END
 END vccd_1p0.gds758
 PIN vccd_1p0.gds759
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.718 17.544 20.778 17.744 ;
 END
 END vccd_1p0.gds759
 PIN vccd_1p0.gds760
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.602 15.7365 24.642 15.9365 ;
 END
 END vccd_1p0.gds760
 PIN vccd_1p0.gds761
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.51 15.778 23.55 15.978 ;
 END
 END vccd_1p0.gds761
 PIN vccd_1p0.gds762
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 18.0025 23.842 18.2025 ;
 END
 END vccd_1p0.gds762
 PIN vccd_1p0.gds763
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 25.004 18.0955 25.06 18.2955 ;
 RECT 24.836 18.0655 24.892 18.2655 ;
 RECT 24.332 18.0955 24.388 18.2955 ;
 RECT 23.996 17.964 24.052 18.164 ;
 RECT 24.164 18.0655 24.22 18.2655 ;
 RECT 24.668 17.964 24.724 18.164 ;
 RECT 23.24 18.0955 23.296 18.2955 ;
 RECT 23.072 18.0655 23.128 18.2655 ;
 RECT 23.576 17.964 23.632 18.164 ;
 RECT 22.568 18.0955 22.624 18.2955 ;
 RECT 22.4 18.0655 22.456 18.2655 ;
 RECT 22.904 17.964 22.96 18.164 ;
 RECT 21.896 18.0955 21.952 18.2955 ;
 RECT 21.728 18.0655 21.784 18.2655 ;
 RECT 22.232 17.964 22.288 18.164 ;
 RECT 21.224 18.0955 21.28 18.2955 ;
 RECT 21.056 18.0655 21.112 18.2655 ;
 RECT 21.56 17.964 21.616 18.164 ;
 RECT 20.552 18.0955 20.608 18.2955 ;
 RECT 20.888 17.964 20.944 18.164 ;
 RECT 20.384 18.0655 20.44 18.2655 ;
 RECT 23.828 17.5945 23.884 17.7945 ;
 END
 END vccd_1p0.gds763
 PIN vccd_1p0.gds764
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.634 15.7365 28.674 15.9365 ;
 END
 END vccd_1p0.gds764
 PIN vccd_1p0.gds765
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.962 15.7365 28.002 15.9365 ;
 END
 END vccd_1p0.gds765
 PIN vccd_1p0.gds766
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.29 15.7365 27.33 15.9365 ;
 END
 END vccd_1p0.gds766
 PIN vccd_1p0.gds767
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.618 15.7365 26.658 15.9365 ;
 END
 END vccd_1p0.gds767
 PIN vccd_1p0.gds768
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.946 15.7365 25.986 15.9365 ;
 END
 END vccd_1p0.gds768
 PIN vccd_1p0.gds769
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.274 15.7365 25.314 15.9365 ;
 END
 END vccd_1p0.gds769
 PIN vccd_1p0.gds770
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.866 17.5755 28.926 17.7755 ;
 END
 END vccd_1p0.gds770
 PIN vccd_1p0.gds771
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.202 17.544 29.262 17.744 ;
 END
 END vccd_1p0.gds771
 PIN vccd_1p0.gds772
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.194 17.5755 28.254 17.7755 ;
 END
 END vccd_1p0.gds772
 PIN vccd_1p0.gds773
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.53 17.544 28.59 17.744 ;
 END
 END vccd_1p0.gds773
 PIN vccd_1p0.gds774
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.522 17.5755 27.582 17.7755 ;
 END
 END vccd_1p0.gds774
 PIN vccd_1p0.gds775
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.858 17.544 27.918 17.744 ;
 END
 END vccd_1p0.gds775
 PIN vccd_1p0.gds776
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.85 17.5755 26.91 17.7755 ;
 END
 END vccd_1p0.gds776
 PIN vccd_1p0.gds777
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.186 17.544 27.246 17.744 ;
 END
 END vccd_1p0.gds777
 PIN vccd_1p0.gds778
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.178 17.5755 26.238 17.7755 ;
 END
 END vccd_1p0.gds778
 PIN vccd_1p0.gds779
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.514 17.544 26.574 17.744 ;
 END
 END vccd_1p0.gds779
 PIN vccd_1p0.gds780
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.506 17.5755 25.566 17.7755 ;
 END
 END vccd_1p0.gds780
 PIN vccd_1p0.gds781
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.842 17.544 25.902 17.744 ;
 END
 END vccd_1p0.gds781
 PIN vccd_1p0.gds782
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 17.3415 29.95 17.5415 ;
 END
 END vccd_1p0.gds782
 PIN vccd_1p0.gds783
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.306 15.7405 29.346 15.9405 ;
 END
 END vccd_1p0.gds783
 PIN vccd_1p0.gds784
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 18.0675 29.706 18.2675 ;
 END
 END vccd_1p0.gds784
 PIN vccd_1p0.gds785
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 29.036 18.0955 29.092 18.2955 ;
 RECT 28.868 18.0655 28.924 18.2655 ;
 RECT 29.372 17.964 29.428 18.164 ;
 RECT 28.364 18.0955 28.42 18.2955 ;
 RECT 28.196 18.0655 28.252 18.2655 ;
 RECT 28.7 17.964 28.756 18.164 ;
 RECT 27.692 18.0955 27.748 18.2955 ;
 RECT 27.524 18.0655 27.58 18.2655 ;
 RECT 28.028 17.964 28.084 18.164 ;
 RECT 27.02 18.0955 27.076 18.2955 ;
 RECT 26.852 18.0655 26.908 18.2655 ;
 RECT 27.356 17.964 27.412 18.164 ;
 RECT 26.348 18.0955 26.404 18.2955 ;
 RECT 26.18 18.0655 26.236 18.2655 ;
 RECT 26.684 17.964 26.74 18.164 ;
 RECT 25.676 18.0955 25.732 18.2955 ;
 RECT 25.508 18.0655 25.564 18.2655 ;
 RECT 26.012 17.964 26.068 18.164 ;
 RECT 25.34 17.964 25.396 18.164 ;
 RECT 30.044 16.967 30.1 17.167 ;
 RECT 29.792 17.5945 29.848 17.7945 ;
 RECT 29.624 17.666 29.68 17.866 ;
 END
 END vccd_1p0.gds785
 PIN vccd_1p0.gds786
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 19.504 31.03 19.704 ;
 END
 END vccd_1p0.gds786
 PIN vccd_1p0.gds787
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 17.697 31.45 17.897 ;
 END
 END vccd_1p0.gds787
 PIN vccd_1p0.gds788
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.386 17.795 33.442 17.995 ;
 END
 END vccd_1p0.gds788
 PIN vccd_1p0.gds789
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 17.1315 33.278 17.3315 ;
 END
 END vccd_1p0.gds789
 PIN vccd_1p0.gds790
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 19.568 33.278 19.768 ;
 END
 END vccd_1p0.gds790
 PIN vccd_1p0.gds791
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 19.504 31.45 19.704 ;
 END
 END vccd_1p0.gds791
 PIN vccd_1p0.gds792
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 18.2 32.794 18.4 ;
 END
 END vccd_1p0.gds792
 PIN vccd_1p0.gds793
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 19.436 32.342 19.636 ;
 END
 END vccd_1p0.gds793
 PIN vccd_1p0.gds794
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 18.5525 30.79 18.7525 ;
 END
 END vccd_1p0.gds794
 PIN vccd_1p0.gds795
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 18.995 30.19 19.195 ;
 END
 END vccd_1p0.gds795
 PIN vccd_1p0.gds796
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 15.453 31.03 15.653 ;
 END
 END vccd_1p0.gds796
 PIN vccd_1p0.gds797
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 18.271 31.03 18.471 ;
 END
 END vccd_1p0.gds797
 PIN vccd_1p0.gds798
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 16.607 31.986 16.807 ;
 END
 END vccd_1p0.gds798
 PIN vccd_1p0.gds799
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 16.7735 31.794 16.9735 ;
 END
 END vccd_1p0.gds799
 PIN vccd_1p0.gds800
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 19.599 35.142 19.799 ;
 END
 END vccd_1p0.gds800
 PIN vccd_1p0.gds801
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 19.4835 35.014 19.6835 ;
 END
 END vccd_1p0.gds801
 PIN vccd_1p0.gds802
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 17.9255 32.55 18.1255 ;
 END
 END vccd_1p0.gds802
 PIN vccd_1p0.gds803
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 19.6315 31.986 19.8315 ;
 END
 END vccd_1p0.gds803
 PIN vccd_1p0.gds804
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 19.232 34.786 19.432 ;
 END
 END vccd_1p0.gds804
 PIN vccd_1p0.gds805
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 17.561 34.626 17.761 ;
 END
 END vccd_1p0.gds805
 PIN vccd_1p0.gds806
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 17.143 34.206 17.343 ;
 END
 END vccd_1p0.gds806
 PIN vccd_1p0.gds807
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 15.8895 35.142 16.0895 ;
 END
 END vccd_1p0.gds807
 PIN vccd_1p0.gds808
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 15.902 35.014 16.102 ;
 END
 END vccd_1p0.gds808
 PIN vccd_1p0.gds809
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 32.312 17.68 32.368 17.88 ;
 RECT 30.296 17.47 30.352 17.67 ;
 RECT 32.144 17.774 32.2 17.974 ;
 RECT 31.976 17.774 32.032 17.974 ;
 RECT 31.808 17.666 31.864 17.866 ;
 RECT 31.64 17.5945 31.696 17.7945 ;
 RECT 31.472 17.5945 31.528 17.7945 ;
 RECT 31.304 17.5945 31.36 17.7945 ;
 RECT 31.136 17.774 31.192 17.974 ;
 RECT 30.968 17.774 31.024 17.974 ;
 RECT 30.8 17.666 30.856 17.866 ;
 RECT 33.824 17.4835 33.88 17.6835 ;
 RECT 33.656 17.4835 33.712 17.6835 ;
 RECT 33.488 17.4835 33.544 17.6835 ;
 RECT 33.32 17.4835 33.376 17.6835 ;
 RECT 33.152 17.4835 33.208 17.6835 ;
 RECT 32.984 17.4835 33.04 17.6835 ;
 RECT 32.816 17.4835 32.872 17.6835 ;
 RECT 32.648 17.5945 32.704 17.7945 ;
 RECT 32.48 17.68 32.536 17.88 ;
 RECT 33.992 17.4835 34.048 17.6835 ;
 RECT 35 17.4975 35.056 17.6975 ;
 RECT 34.832 17.68 34.888 17.88 ;
 RECT 34.664 17.5945 34.72 17.7945 ;
 RECT 34.496 17.5945 34.552 17.7945 ;
 RECT 34.328 17.68 34.384 17.88 ;
 RECT 34.16 17.68 34.216 17.88 ;
 END
 END vccd_1p0.gds809
 PIN vccd_1p0.gds810
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.89 15.7365 39.93 15.9365 ;
 END
 END vccd_1p0.gds810
 PIN vccd_1p0.gds811
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.218 15.7365 39.258 15.9365 ;
 END
 END vccd_1p0.gds811
 PIN vccd_1p0.gds812
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.546 15.7365 38.586 15.9365 ;
 END
 END vccd_1p0.gds812
 PIN vccd_1p0.gds813
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.874 15.7365 37.914 15.9365 ;
 END
 END vccd_1p0.gds813
 PIN vccd_1p0.gds814
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.202 15.7365 37.242 15.9365 ;
 END
 END vccd_1p0.gds814
 PIN vccd_1p0.gds815
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.53 15.7365 36.57 15.9365 ;
 END
 END vccd_1p0.gds815
 PIN vccd_1p0.gds816
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.122 17.5755 40.182 17.7755 ;
 END
 END vccd_1p0.gds816
 PIN vccd_1p0.gds817
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.45 17.5755 39.51 17.7755 ;
 END
 END vccd_1p0.gds817
 PIN vccd_1p0.gds818
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.786 17.544 39.846 17.744 ;
 END
 END vccd_1p0.gds818
 PIN vccd_1p0.gds819
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.778 17.5755 38.838 17.7755 ;
 END
 END vccd_1p0.gds819
 PIN vccd_1p0.gds820
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.114 17.544 39.174 17.744 ;
 END
 END vccd_1p0.gds820
 PIN vccd_1p0.gds821
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.106 17.5755 38.166 17.7755 ;
 END
 END vccd_1p0.gds821
 PIN vccd_1p0.gds822
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.442 17.544 38.502 17.744 ;
 END
 END vccd_1p0.gds822
 PIN vccd_1p0.gds823
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.434 17.5755 37.494 17.7755 ;
 END
 END vccd_1p0.gds823
 PIN vccd_1p0.gds824
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.77 17.544 37.83 17.744 ;
 END
 END vccd_1p0.gds824
 PIN vccd_1p0.gds825
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.762 17.5755 36.822 17.7755 ;
 END
 END vccd_1p0.gds825
 PIN vccd_1p0.gds826
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.098 17.544 37.158 17.744 ;
 END
 END vccd_1p0.gds826
 PIN vccd_1p0.gds827
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.09 17.5755 36.15 17.7755 ;
 END
 END vccd_1p0.gds827
 PIN vccd_1p0.gds828
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.426 17.544 36.486 17.744 ;
 END
 END vccd_1p0.gds828
 PIN vccd_1p0.gds829
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.418 17.4515 35.478 17.6515 ;
 END
 END vccd_1p0.gds829
 PIN vccd_1p0.gds830
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.754 17.544 35.814 17.744 ;
 END
 END vccd_1p0.gds830
 PIN vccd_1p0.gds831
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.858 15.7365 35.898 15.9365 ;
 END
 END vccd_1p0.gds831
 PIN vccd_1p0.gds832
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 40.124 18.0655 40.18 18.2655 ;
 RECT 39.62 18.0955 39.676 18.2955 ;
 RECT 39.452 18.0655 39.508 18.2655 ;
 RECT 39.956 17.964 40.012 18.164 ;
 RECT 38.948 18.0955 39.004 18.2955 ;
 RECT 38.78 18.0655 38.836 18.2655 ;
 RECT 39.284 17.964 39.34 18.164 ;
 RECT 38.276 18.0955 38.332 18.2955 ;
 RECT 38.108 18.0655 38.164 18.2655 ;
 RECT 38.612 17.964 38.668 18.164 ;
 RECT 37.604 18.0955 37.66 18.2955 ;
 RECT 37.436 18.0655 37.492 18.2655 ;
 RECT 37.94 17.964 37.996 18.164 ;
 RECT 36.932 18.0955 36.988 18.2955 ;
 RECT 36.764 18.0655 36.82 18.2655 ;
 RECT 37.268 17.964 37.324 18.164 ;
 RECT 36.26 18.0955 36.316 18.2955 ;
 RECT 36.092 18.0655 36.148 18.2655 ;
 RECT 36.596 17.964 36.652 18.164 ;
 RECT 35.588 18.0955 35.644 18.2955 ;
 RECT 35.252 17.964 35.308 18.164 ;
 RECT 35.42 18.0655 35.476 18.2655 ;
 RECT 35.924 17.964 35.98 18.164 ;
 END
 END vccd_1p0.gds832
 PIN vccd_1p0.gds833
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.014 15.7365 45.054 15.9365 ;
 END
 END vccd_1p0.gds833
 PIN vccd_1p0.gds834
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.342 15.7365 44.382 15.9365 ;
 END
 END vccd_1p0.gds834
 PIN vccd_1p0.gds835
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.67 15.7365 43.71 15.9365 ;
 END
 END vccd_1p0.gds835
 PIN vccd_1p0.gds836
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.998 15.7365 43.038 15.9365 ;
 END
 END vccd_1p0.gds836
 PIN vccd_1p0.gds837
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.326 15.7365 42.366 15.9365 ;
 END
 END vccd_1p0.gds837
 PIN vccd_1p0.gds838
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.574 17.5755 44.634 17.7755 ;
 END
 END vccd_1p0.gds838
 PIN vccd_1p0.gds839
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.91 17.544 44.97 17.744 ;
 END
 END vccd_1p0.gds839
 PIN vccd_1p0.gds840
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.902 17.5755 43.962 17.7755 ;
 END
 END vccd_1p0.gds840
 PIN vccd_1p0.gds841
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.238 17.544 44.298 17.744 ;
 END
 END vccd_1p0.gds841
 PIN vccd_1p0.gds842
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.23 17.5755 43.29 17.7755 ;
 END
 END vccd_1p0.gds842
 PIN vccd_1p0.gds843
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.566 17.544 43.626 17.744 ;
 END
 END vccd_1p0.gds843
 PIN vccd_1p0.gds844
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.558 17.5755 42.618 17.7755 ;
 END
 END vccd_1p0.gds844
 PIN vccd_1p0.gds845
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.894 17.544 42.954 17.744 ;
 END
 END vccd_1p0.gds845
 PIN vccd_1p0.gds846
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.886 17.5755 41.946 17.7755 ;
 END
 END vccd_1p0.gds846
 PIN vccd_1p0.gds847
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.222 17.544 42.282 17.744 ;
 END
 END vccd_1p0.gds847
 PIN vccd_1p0.gds848
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.214 17.5755 41.274 17.7755 ;
 END
 END vccd_1p0.gds848
 PIN vccd_1p0.gds849
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.55 17.544 41.61 17.744 ;
 END
 END vccd_1p0.gds849
 PIN vccd_1p0.gds850
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.458 17.544 40.518 17.744 ;
 END
 END vccd_1p0.gds850
 PIN vccd_1p0.gds851
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 18.0025 40.894 18.2025 ;
 END
 END vccd_1p0.gds851
 PIN vccd_1p0.gds852
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.654 15.7365 41.694 15.9365 ;
 END
 END vccd_1p0.gds852
 PIN vccd_1p0.gds853
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.562 15.778 40.602 15.978 ;
 END
 END vccd_1p0.gds853
 PIN vccd_1p0.gds854
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 44.744 18.0955 44.8 18.2955 ;
 RECT 44.576 18.0655 44.632 18.2655 ;
 RECT 45.08 17.964 45.136 18.164 ;
 RECT 44.072 18.0955 44.128 18.2955 ;
 RECT 43.904 18.0655 43.96 18.2655 ;
 RECT 44.408 17.964 44.464 18.164 ;
 RECT 43.4 18.0955 43.456 18.2955 ;
 RECT 43.232 18.0655 43.288 18.2655 ;
 RECT 43.736 17.964 43.792 18.164 ;
 RECT 42.728 18.0955 42.784 18.2955 ;
 RECT 42.56 18.0655 42.616 18.2655 ;
 RECT 43.064 17.964 43.12 18.164 ;
 RECT 42.056 18.0955 42.112 18.2955 ;
 RECT 41.888 18.0655 41.944 18.2655 ;
 RECT 42.392 17.964 42.448 18.164 ;
 RECT 41.384 18.0955 41.44 18.2955 ;
 RECT 41.048 17.964 41.104 18.164 ;
 RECT 41.216 18.0655 41.272 18.2655 ;
 RECT 41.72 17.964 41.776 18.164 ;
 RECT 40.628 17.964 40.684 18.164 ;
 RECT 40.292 18.0955 40.348 18.2955 ;
 RECT 40.88 17.5945 40.936 17.7945 ;
 END
 END vccd_1p0.gds854
 PIN vccd_1p0.gds855
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.686 15.7365 45.726 15.9365 ;
 END
 END vccd_1p0.gds855
 PIN vccd_1p0.gds856
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.918 17.5755 45.978 17.7755 ;
 END
 END vccd_1p0.gds856
 PIN vccd_1p0.gds857
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.254 17.544 46.314 17.744 ;
 END
 END vccd_1p0.gds857
 PIN vccd_1p0.gds858
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.246 17.5755 45.306 17.7755 ;
 END
 END vccd_1p0.gds858
 PIN vccd_1p0.gds859
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.582 17.544 45.642 17.744 ;
 END
 END vccd_1p0.gds859
 PIN vccd_1p0.gds860
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 17.697 48.502 17.897 ;
 END
 END vccd_1p0.gds860
 PIN vccd_1p0.gds861
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 19.504 48.082 19.704 ;
 END
 END vccd_1p0.gds861
 PIN vccd_1p0.gds862
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 19.504 48.502 19.704 ;
 END
 END vccd_1p0.gds862
 PIN vccd_1p0.gds863
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 18.2 49.846 18.4 ;
 END
 END vccd_1p0.gds863
 PIN vccd_1p0.gds864
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 19.436 49.394 19.636 ;
 END
 END vccd_1p0.gds864
 PIN vccd_1p0.gds865
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 18.5525 47.842 18.7525 ;
 END
 END vccd_1p0.gds865
 PIN vccd_1p0.gds866
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 18.995 47.242 19.195 ;
 END
 END vccd_1p0.gds866
 PIN vccd_1p0.gds867
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 17.3415 47.002 17.5415 ;
 END
 END vccd_1p0.gds867
 PIN vccd_1p0.gds868
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 15.453 48.082 15.653 ;
 END
 END vccd_1p0.gds868
 PIN vccd_1p0.gds869
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 18.271 48.082 18.471 ;
 END
 END vccd_1p0.gds869
 PIN vccd_1p0.gds870
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 16.607 49.038 16.807 ;
 END
 END vccd_1p0.gds870
 PIN vccd_1p0.gds871
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.358 15.7405 46.398 15.9405 ;
 END
 END vccd_1p0.gds871
 PIN vccd_1p0.gds872
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 16.7735 48.846 16.9735 ;
 END
 END vccd_1p0.gds872
 PIN vccd_1p0.gds873
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 19.6315 49.038 19.8315 ;
 END
 END vccd_1p0.gds873
 PIN vccd_1p0.gds874
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 17.9255 49.602 18.1255 ;
 END
 END vccd_1p0.gds874
 PIN vccd_1p0.gds875
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 18.0675 46.758 18.2675 ;
 END
 END vccd_1p0.gds875
 PIN vccd_1p0.gds876
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 17.1315 50.33 17.3315 ;
 END
 END vccd_1p0.gds876
 PIN vccd_1p0.gds877
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 46.088 18.0955 46.144 18.2955 ;
 RECT 45.92 18.0655 45.976 18.2655 ;
 RECT 46.424 17.964 46.48 18.164 ;
 RECT 45.416 18.0955 45.472 18.2955 ;
 RECT 45.248 18.0655 45.304 18.2655 ;
 RECT 45.752 17.964 45.808 18.164 ;
 RECT 47.096 16.967 47.152 17.167 ;
 RECT 49.364 17.68 49.42 17.88 ;
 RECT 46.844 17.5945 46.9 17.7945 ;
 RECT 47.348 17.47 47.404 17.67 ;
 RECT 46.676 17.666 46.732 17.866 ;
 RECT 49.196 17.774 49.252 17.974 ;
 RECT 49.028 17.774 49.084 17.974 ;
 RECT 48.86 17.666 48.916 17.866 ;
 RECT 48.692 17.5945 48.748 17.7945 ;
 RECT 48.524 17.5945 48.58 17.7945 ;
 RECT 48.356 17.5945 48.412 17.7945 ;
 RECT 48.188 17.774 48.244 17.974 ;
 RECT 48.02 17.774 48.076 17.974 ;
 RECT 47.852 17.666 47.908 17.866 ;
 RECT 50.204 17.4835 50.26 17.6835 ;
 RECT 50.036 17.4835 50.092 17.6835 ;
 RECT 49.868 17.4835 49.924 17.6835 ;
 RECT 49.7 17.5945 49.756 17.7945 ;
 RECT 49.532 17.68 49.588 17.88 ;
 END
 END vccd_1p0.gds877
 PIN vccd_1p0.gds878
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.926 15.7365 54.966 15.9365 ;
 END
 END vccd_1p0.gds878
 PIN vccd_1p0.gds879
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.254 15.7365 54.294 15.9365 ;
 END
 END vccd_1p0.gds879
 PIN vccd_1p0.gds880
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.582 15.7365 53.622 15.9365 ;
 END
 END vccd_1p0.gds880
 PIN vccd_1p0.gds881
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.158 17.5755 55.218 17.7755 ;
 END
 END vccd_1p0.gds881
 PIN vccd_1p0.gds882
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.486 17.5755 54.546 17.7755 ;
 END
 END vccd_1p0.gds882
 PIN vccd_1p0.gds883
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.822 17.544 54.882 17.744 ;
 END
 END vccd_1p0.gds883
 PIN vccd_1p0.gds884
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.814 17.5755 53.874 17.7755 ;
 END
 END vccd_1p0.gds884
 PIN vccd_1p0.gds885
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.15 17.544 54.21 17.744 ;
 END
 END vccd_1p0.gds885
 PIN vccd_1p0.gds886
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.142 17.5755 53.202 17.7755 ;
 END
 END vccd_1p0.gds886
 PIN vccd_1p0.gds887
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.478 17.544 53.538 17.744 ;
 END
 END vccd_1p0.gds887
 PIN vccd_1p0.gds888
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.47 17.4515 52.53 17.6515 ;
 END
 END vccd_1p0.gds888
 PIN vccd_1p0.gds889
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.806 17.544 52.866 17.744 ;
 END
 END vccd_1p0.gds889
 PIN vccd_1p0.gds890
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.438 17.795 50.494 17.995 ;
 END
 END vccd_1p0.gds890
 PIN vccd_1p0.gds891
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 19.568 50.33 19.768 ;
 END
 END vccd_1p0.gds891
 PIN vccd_1p0.gds892
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 15.8895 52.194 16.0895 ;
 END
 END vccd_1p0.gds892
 PIN vccd_1p0.gds893
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 15.902 52.066 16.102 ;
 END
 END vccd_1p0.gds893
 PIN vccd_1p0.gds894
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 17.4875 51.678 17.6875 ;
 END
 END vccd_1p0.gds894
 PIN vccd_1p0.gds895
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 19.599 52.194 19.799 ;
 END
 END vccd_1p0.gds895
 PIN vccd_1p0.gds896
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 19.4835 52.066 19.6835 ;
 END
 END vccd_1p0.gds896
 PIN vccd_1p0.gds897
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 17.143 51.258 17.343 ;
 END
 END vccd_1p0.gds897
 PIN vccd_1p0.gds898
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 19.3655 51.838 19.5655 ;
 END
 END vccd_1p0.gds898
 PIN vccd_1p0.gds899
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.91 15.7365 52.95 15.9365 ;
 END
 END vccd_1p0.gds899
 PIN vccd_1p0.gds900
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 55.16 18.0655 55.216 18.2655 ;
 RECT 54.656 18.0955 54.712 18.2955 ;
 RECT 54.488 18.0655 54.544 18.2655 ;
 RECT 54.992 17.964 55.048 18.164 ;
 RECT 53.984 18.0955 54.04 18.2955 ;
 RECT 53.816 18.0655 53.872 18.2655 ;
 RECT 54.32 17.964 54.376 18.164 ;
 RECT 53.312 18.0955 53.368 18.2955 ;
 RECT 53.144 18.0655 53.2 18.2655 ;
 RECT 53.648 17.964 53.704 18.164 ;
 RECT 52.64 18.0955 52.696 18.2955 ;
 RECT 52.304 17.964 52.36 18.164 ;
 RECT 52.472 18.0655 52.528 18.2655 ;
 RECT 52.976 17.964 53.032 18.164 ;
 RECT 50.876 17.4835 50.932 17.6835 ;
 RECT 50.708 17.4835 50.764 17.6835 ;
 RECT 50.54 17.4835 50.596 17.6835 ;
 RECT 50.372 17.4835 50.428 17.6835 ;
 RECT 51.044 17.4835 51.1 17.6835 ;
 RECT 52.052 17.4975 52.108 17.6975 ;
 RECT 51.884 17.68 51.94 17.88 ;
 RECT 51.716 17.5945 51.772 17.7945 ;
 RECT 51.548 17.5945 51.604 17.7945 ;
 RECT 51.38 17.68 51.436 17.88 ;
 RECT 51.212 17.68 51.268 17.88 ;
 END
 END vccd_1p0.gds900
 PIN vccd_1p0.gds901
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.05 15.7365 60.09 15.9365 ;
 END
 END vccd_1p0.gds901
 PIN vccd_1p0.gds902
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.378 15.7365 59.418 15.9365 ;
 END
 END vccd_1p0.gds902
 PIN vccd_1p0.gds903
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.942 15.7365 56.982 15.9365 ;
 END
 END vccd_1p0.gds903
 PIN vccd_1p0.gds904
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.27 15.7365 56.31 15.9365 ;
 END
 END vccd_1p0.gds904
 PIN vccd_1p0.gds905
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.598 15.7365 55.638 15.9365 ;
 END
 END vccd_1p0.gds905
 PIN vccd_1p0.gds906
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.61 17.5755 59.67 17.7755 ;
 END
 END vccd_1p0.gds906
 PIN vccd_1p0.gds907
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.946 17.544 60.006 17.744 ;
 END
 END vccd_1p0.gds907
 PIN vccd_1p0.gds908
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.938 17.5755 58.998 17.7755 ;
 END
 END vccd_1p0.gds908
 PIN vccd_1p0.gds909
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.274 17.544 59.334 17.744 ;
 END
 END vccd_1p0.gds909
 PIN vccd_1p0.gds910
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.266 17.5755 58.326 17.7755 ;
 END
 END vccd_1p0.gds910
 PIN vccd_1p0.gds911
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.602 17.544 58.662 17.744 ;
 END
 END vccd_1p0.gds911
 PIN vccd_1p0.gds912
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.174 17.5755 57.234 17.7755 ;
 END
 END vccd_1p0.gds912
 PIN vccd_1p0.gds913
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.51 17.544 57.57 17.744 ;
 END
 END vccd_1p0.gds913
 PIN vccd_1p0.gds914
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.502 17.5755 56.562 17.7755 ;
 END
 END vccd_1p0.gds914
 PIN vccd_1p0.gds915
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.838 17.544 56.898 17.744 ;
 END
 END vccd_1p0.gds915
 PIN vccd_1p0.gds916
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.83 17.5755 55.89 17.7755 ;
 END
 END vccd_1p0.gds916
 PIN vccd_1p0.gds917
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.166 17.544 56.226 17.744 ;
 END
 END vccd_1p0.gds917
 PIN vccd_1p0.gds918
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.494 17.544 55.554 17.744 ;
 END
 END vccd_1p0.gds918
 PIN vccd_1p0.gds919
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.706 15.7365 58.746 15.9365 ;
 END
 END vccd_1p0.gds919
 PIN vccd_1p0.gds920
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.614 15.778 57.654 15.978 ;
 END
 END vccd_1p0.gds920
 PIN vccd_1p0.gds921
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 18.0025 57.946 18.2025 ;
 END
 END vccd_1p0.gds921
 PIN vccd_1p0.gds922
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 59.78 18.0955 59.836 18.2955 ;
 RECT 59.612 18.0655 59.668 18.2655 ;
 RECT 60.116 17.964 60.172 18.164 ;
 RECT 59.108 18.0955 59.164 18.2955 ;
 RECT 58.94 18.0655 58.996 18.2655 ;
 RECT 59.444 17.964 59.5 18.164 ;
 RECT 58.436 18.0955 58.492 18.2955 ;
 RECT 58.1 17.964 58.156 18.164 ;
 RECT 58.268 18.0655 58.324 18.2655 ;
 RECT 58.772 17.964 58.828 18.164 ;
 RECT 57.344 18.0955 57.4 18.2955 ;
 RECT 57.176 18.0655 57.232 18.2655 ;
 RECT 57.68 17.964 57.736 18.164 ;
 RECT 56.672 18.0955 56.728 18.2955 ;
 RECT 56.504 18.0655 56.56 18.2655 ;
 RECT 57.008 17.964 57.064 18.164 ;
 RECT 56 18.0955 56.056 18.2955 ;
 RECT 55.832 18.0655 55.888 18.2655 ;
 RECT 56.336 17.964 56.392 18.164 ;
 RECT 55.328 18.0955 55.384 18.2955 ;
 RECT 55.664 17.964 55.72 18.164 ;
 RECT 57.932 17.5945 57.988 17.7945 ;
 END
 END vccd_1p0.gds922
 PIN vccd_1p0.gds923
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.738 15.7365 62.778 15.9365 ;
 END
 END vccd_1p0.gds923
 PIN vccd_1p0.gds924
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.066 15.7365 62.106 15.9365 ;
 END
 END vccd_1p0.gds924
 PIN vccd_1p0.gds925
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.394 15.7365 61.434 15.9365 ;
 END
 END vccd_1p0.gds925
 PIN vccd_1p0.gds926
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.722 15.7365 60.762 15.9365 ;
 END
 END vccd_1p0.gds926
 PIN vccd_1p0.gds927
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.97 17.5755 63.03 17.7755 ;
 END
 END vccd_1p0.gds927
 PIN vccd_1p0.gds928
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.306 17.544 63.366 17.744 ;
 END
 END vccd_1p0.gds928
 PIN vccd_1p0.gds929
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.298 17.5755 62.358 17.7755 ;
 END
 END vccd_1p0.gds929
 PIN vccd_1p0.gds930
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.634 17.544 62.694 17.744 ;
 END
 END vccd_1p0.gds930
 PIN vccd_1p0.gds931
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.626 17.5755 61.686 17.7755 ;
 END
 END vccd_1p0.gds931
 PIN vccd_1p0.gds932
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.962 17.544 62.022 17.744 ;
 END
 END vccd_1p0.gds932
 PIN vccd_1p0.gds933
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.954 17.5755 61.014 17.7755 ;
 END
 END vccd_1p0.gds933
 PIN vccd_1p0.gds934
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.29 17.544 61.35 17.744 ;
 END
 END vccd_1p0.gds934
 PIN vccd_1p0.gds935
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.282 17.5755 60.342 17.7755 ;
 END
 END vccd_1p0.gds935
 PIN vccd_1p0.gds936
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.618 17.544 60.678 17.744 ;
 END
 END vccd_1p0.gds936
 PIN vccd_1p0.gds937
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 19.504 65.134 19.704 ;
 END
 END vccd_1p0.gds937
 PIN vccd_1p0.gds938
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 18.5525 64.894 18.7525 ;
 END
 END vccd_1p0.gds938
 PIN vccd_1p0.gds939
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 18.995 64.294 19.195 ;
 END
 END vccd_1p0.gds939
 PIN vccd_1p0.gds940
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 18.0675 63.81 18.2675 ;
 END
 END vccd_1p0.gds940
 PIN vccd_1p0.gds941
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 17.3415 64.054 17.5415 ;
 END
 END vccd_1p0.gds941
 PIN vccd_1p0.gds942
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 15.453 65.134 15.653 ;
 END
 END vccd_1p0.gds942
 PIN vccd_1p0.gds943
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 18.271 65.134 18.471 ;
 END
 END vccd_1p0.gds943
 PIN vccd_1p0.gds944
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.41 15.7405 63.45 15.9405 ;
 END
 END vccd_1p0.gds944
 PIN vccd_1p0.gds945
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 63.14 18.0955 63.196 18.2955 ;
 RECT 62.972 18.0655 63.028 18.2655 ;
 RECT 63.476 17.964 63.532 18.164 ;
 RECT 62.468 18.0955 62.524 18.2955 ;
 RECT 62.3 18.0655 62.356 18.2655 ;
 RECT 62.804 17.964 62.86 18.164 ;
 RECT 61.796 18.0955 61.852 18.2955 ;
 RECT 61.628 18.0655 61.684 18.2655 ;
 RECT 62.132 17.964 62.188 18.164 ;
 RECT 61.124 18.0955 61.18 18.2955 ;
 RECT 60.956 18.0655 61.012 18.2655 ;
 RECT 61.46 17.964 61.516 18.164 ;
 RECT 60.452 18.0955 60.508 18.2955 ;
 RECT 60.788 17.964 60.844 18.164 ;
 RECT 60.284 18.0655 60.34 18.2655 ;
 RECT 64.148 16.967 64.204 17.167 ;
 RECT 63.896 17.5945 63.952 17.7945 ;
 RECT 64.4 17.47 64.456 17.67 ;
 RECT 63.728 17.666 63.784 17.866 ;
 RECT 65.072 17.774 65.128 17.974 ;
 RECT 64.904 17.666 64.96 17.866 ;
 END
 END vccd_1p0.gds945
 PIN vccd_1p0.gds946
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.194 17.5755 70.254 17.7755 ;
 END
 END vccd_1p0.gds946
 PIN vccd_1p0.gds947
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.522 17.4515 69.582 17.6515 ;
 END
 END vccd_1p0.gds947
 PIN vccd_1p0.gds948
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.858 17.544 69.918 17.744 ;
 END
 END vccd_1p0.gds948
 PIN vccd_1p0.gds949
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 15.8895 69.246 16.0895 ;
 END
 END vccd_1p0.gds949
 PIN vccd_1p0.gds950
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 15.902 69.118 16.102 ;
 END
 END vccd_1p0.gds950
 PIN vccd_1p0.gds951
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 17.697 65.554 17.897 ;
 END
 END vccd_1p0.gds951
 PIN vccd_1p0.gds952
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 19.568 67.382 19.768 ;
 END
 END vccd_1p0.gds952
 PIN vccd_1p0.gds953
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 19.504 65.554 19.704 ;
 END
 END vccd_1p0.gds953
 PIN vccd_1p0.gds954
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 19.436 66.446 19.636 ;
 END
 END vccd_1p0.gds954
 PIN vccd_1p0.gds955
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 16.607 66.09 16.807 ;
 END
 END vccd_1p0.gds955
 PIN vccd_1p0.gds956
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 16.7735 65.898 16.9735 ;
 END
 END vccd_1p0.gds956
 PIN vccd_1p0.gds957
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 17.4875 68.73 17.6875 ;
 END
 END vccd_1p0.gds957
 PIN vccd_1p0.gds958
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 19.599 69.246 19.799 ;
 END
 END vccd_1p0.gds958
 PIN vccd_1p0.gds959
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 19.4835 69.118 19.6835 ;
 END
 END vccd_1p0.gds959
 PIN vccd_1p0.gds960
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 17.143 68.31 17.343 ;
 END
 END vccd_1p0.gds960
 PIN vccd_1p0.gds961
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 17.9255 66.654 18.1255 ;
 END
 END vccd_1p0.gds961
 PIN vccd_1p0.gds962
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 19.6315 66.09 19.8315 ;
 END
 END vccd_1p0.gds962
 PIN vccd_1p0.gds963
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 19.3655 68.89 19.5655 ;
 END
 END vccd_1p0.gds963
 PIN vccd_1p0.gds964
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 18.2 66.898 18.4 ;
 END
 END vccd_1p0.gds964
 PIN vccd_1p0.gds965
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.49 17.795 67.546 17.995 ;
 END
 END vccd_1p0.gds965
 PIN vccd_1p0.gds966
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 17.1315 67.382 17.3315 ;
 END
 END vccd_1p0.gds966
 PIN vccd_1p0.gds967
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.962 15.7365 70.002 15.9365 ;
 END
 END vccd_1p0.gds967
 PIN vccd_1p0.gds968
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 70.196 18.0655 70.252 18.2655 ;
 RECT 69.692 18.0955 69.748 18.2955 ;
 RECT 69.356 17.964 69.412 18.164 ;
 RECT 69.524 18.0655 69.58 18.2655 ;
 RECT 70.028 17.964 70.084 18.164 ;
 RECT 66.416 17.68 66.472 17.88 ;
 RECT 66.248 17.774 66.304 17.974 ;
 RECT 66.08 17.774 66.136 17.974 ;
 RECT 65.912 17.666 65.968 17.866 ;
 RECT 65.744 17.5945 65.8 17.7945 ;
 RECT 65.576 17.5945 65.632 17.7945 ;
 RECT 65.408 17.5945 65.464 17.7945 ;
 RECT 65.24 17.774 65.296 17.974 ;
 RECT 67.928 17.4835 67.984 17.6835 ;
 RECT 67.76 17.4835 67.816 17.6835 ;
 RECT 67.592 17.4835 67.648 17.6835 ;
 RECT 67.424 17.4835 67.48 17.6835 ;
 RECT 67.256 17.4835 67.312 17.6835 ;
 RECT 67.088 17.4835 67.144 17.6835 ;
 RECT 66.92 17.4835 66.976 17.6835 ;
 RECT 66.752 17.5945 66.808 17.7945 ;
 RECT 66.584 17.68 66.64 17.88 ;
 RECT 68.096 17.4835 68.152 17.6835 ;
 RECT 69.104 17.4975 69.16 17.6975 ;
 RECT 68.936 17.68 68.992 17.88 ;
 RECT 68.768 17.5945 68.824 17.7945 ;
 RECT 68.6 17.5945 68.656 17.7945 ;
 RECT 68.432 17.68 68.488 17.88 ;
 RECT 68.264 17.68 68.32 17.88 ;
 END
 END vccd_1p0.gds968
 PIN vccd_1p0.gds969
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.666 15.778 74.706 15.978 ;
 END
 END vccd_1p0.gds969
 PIN vccd_1p0.gds970
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.994 15.7365 74.034 15.9365 ;
 END
 END vccd_1p0.gds970
 PIN vccd_1p0.gds971
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.322 15.7365 73.362 15.9365 ;
 END
 END vccd_1p0.gds971
 PIN vccd_1p0.gds972
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.65 15.7365 72.69 15.9365 ;
 END
 END vccd_1p0.gds972
 PIN vccd_1p0.gds973
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.978 15.7365 72.018 15.9365 ;
 END
 END vccd_1p0.gds973
 PIN vccd_1p0.gds974
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.306 15.7365 71.346 15.9365 ;
 END
 END vccd_1p0.gds974
 PIN vccd_1p0.gds975
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.634 15.7365 70.674 15.9365 ;
 END
 END vccd_1p0.gds975
 PIN vccd_1p0.gds976
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.226 17.5755 74.286 17.7755 ;
 END
 END vccd_1p0.gds976
 PIN vccd_1p0.gds977
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.562 17.544 74.622 17.744 ;
 END
 END vccd_1p0.gds977
 PIN vccd_1p0.gds978
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.554 17.5755 73.614 17.7755 ;
 END
 END vccd_1p0.gds978
 PIN vccd_1p0.gds979
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.89 17.544 73.95 17.744 ;
 END
 END vccd_1p0.gds979
 PIN vccd_1p0.gds980
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.882 17.5755 72.942 17.7755 ;
 END
 END vccd_1p0.gds980
 PIN vccd_1p0.gds981
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.218 17.544 73.278 17.744 ;
 END
 END vccd_1p0.gds981
 PIN vccd_1p0.gds982
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.21 17.5755 72.27 17.7755 ;
 END
 END vccd_1p0.gds982
 PIN vccd_1p0.gds983
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.546 17.544 72.606 17.744 ;
 END
 END vccd_1p0.gds983
 PIN vccd_1p0.gds984
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.538 17.5755 71.598 17.7755 ;
 END
 END vccd_1p0.gds984
 PIN vccd_1p0.gds985
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.874 17.544 71.934 17.744 ;
 END
 END vccd_1p0.gds985
 PIN vccd_1p0.gds986
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.866 17.5755 70.926 17.7755 ;
 END
 END vccd_1p0.gds986
 PIN vccd_1p0.gds987
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.202 17.544 71.262 17.744 ;
 END
 END vccd_1p0.gds987
 PIN vccd_1p0.gds988
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.53 17.544 70.59 17.744 ;
 END
 END vccd_1p0.gds988
 PIN vccd_1p0.gds989
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 74.396 18.0955 74.452 18.2955 ;
 RECT 74.228 18.0655 74.284 18.2655 ;
 RECT 74.732 17.964 74.788 18.164 ;
 RECT 73.724 18.0955 73.78 18.2955 ;
 RECT 73.556 18.0655 73.612 18.2655 ;
 RECT 74.06 17.964 74.116 18.164 ;
 RECT 73.052 18.0955 73.108 18.2955 ;
 RECT 72.884 18.0655 72.94 18.2655 ;
 RECT 73.388 17.964 73.444 18.164 ;
 RECT 72.38 18.0955 72.436 18.2955 ;
 RECT 72.212 18.0655 72.268 18.2655 ;
 RECT 72.716 17.964 72.772 18.164 ;
 RECT 71.708 18.0955 71.764 18.2955 ;
 RECT 71.54 18.0655 71.596 18.2655 ;
 RECT 72.044 17.964 72.1 18.164 ;
 RECT 71.036 18.0955 71.092 18.2955 ;
 RECT 70.868 18.0655 70.924 18.2655 ;
 RECT 71.372 17.964 71.428 18.164 ;
 RECT 70.364 18.0955 70.42 18.2955 ;
 RECT 70.7 17.964 70.756 18.164 ;
 END
 END vccd_1p0.gds989
 PIN vccd_1p0.gds990
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 23.138 0.43 23.338 ;
 END
 END vccd_1p0.gds990
 PIN vccd_1p0.gds991
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 22.937 1.542 23.137 ;
 END
 END vccd_1p0.gds991
 PIN vccd_1p0.gds992
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 23.438 0.548 23.638 ;
 END
 END vccd_1p0.gds992
 PIN vccd_1p0.gds993
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 21.677 1.542 21.877 ;
 END
 END vccd_1p0.gds993
 PIN vccd_1p0.gds994
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 21.5595 5.202 21.7595 ;
 END
 END vccd_1p0.gds994
 PIN vccd_1p0.gds995
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 24.197 1.542 24.397 ;
 END
 END vccd_1p0.gds995
 PIN vccd_1p0.gds996
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 24.0795 5.202 24.2795 ;
 END
 END vccd_1p0.gds996
 PIN vccd_1p0.gds997
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 23.0845 0.858 23.2845 ;
 END
 END vccd_1p0.gds997
 PIN vccd_1p0.gds998
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 23.132 1.362 23.332 ;
 END
 END vccd_1p0.gds998
 PIN vccd_1p0.gds999
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 23.021 1.218 23.221 ;
 END
 END vccd_1p0.gds999
 PIN vccd_1p0.gds1000
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 23.098 1.09 23.298 ;
 END
 END vccd_1p0.gds1000
 PIN vccd_1p0.gds1001
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 24.526 1.782 24.726 ;
 END
 END vccd_1p0.gds1001
 PIN vccd_1p0.gds1002
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 22.8195 5.202 23.0195 ;
 END
 END vccd_1p0.gds1002
 PIN vccd_1p0.gds1003
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 25.1445 2.202 25.3445 ;
 END
 END vccd_1p0.gds1003
 PIN vccd_1p0.gds1004
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 22.869 2.622 23.069 ;
 END
 END vccd_1p0.gds1004
 PIN vccd_1p0.gds1005
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 25.3395 5.202 25.5395 ;
 END
 END vccd_1p0.gds1005
 PIN vccd_1p0.gds1006
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 20.9905 3.666 21.1905 ;
 END
 END vccd_1p0.gds1006
 PIN vccd_1p0.gds1007
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 21.011 4.738 21.211 ;
 END
 END vccd_1p0.gds1007
 PIN vccd_1p0.gds1008
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 25.3585 2.462 25.5585 ;
 END
 END vccd_1p0.gds1008
 PIN vccd_1p0.gds1009
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 22.591 1.962 22.791 ;
 END
 END vccd_1p0.gds1009
 PIN vccd_1p0.gds1010
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 22.9255 3.042 23.1255 ;
 END
 END vccd_1p0.gds1010
 PIN vccd_1p0.gds1011
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 22.928 2.882 23.128 ;
 END
 END vccd_1p0.gds1011
 PIN vccd_1p0.gds1012
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 23.05 3.262 23.25 ;
 END
 END vccd_1p0.gds1012
 PIN vccd_1p0.gds1013
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 23.014 3.39 23.214 ;
 END
 END vccd_1p0.gds1013
 PIN vccd_1p0.gds1014
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 23.0165 3.858 23.2165 ;
 END
 END vccd_1p0.gds1014
 PIN vccd_1p0.gds1015
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 21.668 4.258 21.868 ;
 END
 END vccd_1p0.gds1015
 PIN vccd_1p0.gds1016
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 20.58 4.066 20.78 ;
 END
 END vccd_1p0.gds1016
 PIN vccd_1p0.gds1017
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 23.022 4.546 23.222 ;
 END
 END vccd_1p0.gds1017
 PIN vccd_1p0.gds1018
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 23.026 5.01 23.226 ;
 END
 END vccd_1p0.gds1018
 PIN vccd_1p0.gds1019
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 4.76 20.5015 4.816 20.7015 ;
 RECT 4.928 20.5015 4.984 20.7015 ;
 RECT 4.34 20.542 4.396 20.742 ;
 RECT 3.584 24.2235 3.64 24.4235 ;
 RECT 3.584 22.9635 3.64 23.1635 ;
 RECT 3.584 21.7035 3.64 21.9035 ;
 RECT 4.34 24.322 4.396 24.522 ;
 RECT 4.172 24.322 4.228 24.522 ;
 RECT 4.76 24.2815 4.816 24.4815 ;
 RECT 5.096 24.322 5.152 24.522 ;
 RECT 4.928 24.2815 4.984 24.4815 ;
 RECT 4.34 23.062 4.396 23.262 ;
 RECT 4.172 23.062 4.228 23.262 ;
 RECT 4.76 23.0215 4.816 23.2215 ;
 RECT 5.096 23.062 5.152 23.262 ;
 RECT 4.928 23.0215 4.984 23.2215 ;
 RECT 4.34 21.802 4.396 22.002 ;
 RECT 4.172 21.802 4.228 22.002 ;
 RECT 4.76 21.7615 4.816 21.9615 ;
 RECT 5.096 21.802 5.152 22.002 ;
 RECT 4.928 21.7615 4.984 21.9615 ;
 RECT 4.172 20.542 4.228 20.742 ;
 RECT 5.096 20.542 5.152 20.742 ;
 END
 END vccd_1p0.gds1019
 PIN vccd_1p0.gds1020
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 23.0165 6.838 23.2165 ;
 END
 END vccd_1p0.gds1020
 PIN vccd_1p0.gds1021
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 25.366 6.05 25.566 ;
 END
 END vccd_1p0.gds1021
 PIN vccd_1p0.gds1022
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.754 21.2165 5.794 21.4165 ;
 END
 END vccd_1p0.gds1022
 PIN vccd_1p0.gds1023
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 20.947 5.41 21.147 ;
 END
 END vccd_1p0.gds1023
 PIN vccd_1p0.gds1024
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 24.944 5.922 25.144 ;
 END
 END vccd_1p0.gds1024
 PIN vccd_1p0.gds1025
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 23.1535 5.602 23.3535 ;
 END
 END vccd_1p0.gds1025
 PIN vccd_1p0.gds1026
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 24.053 6.306 24.253 ;
 END
 END vccd_1p0.gds1026
 PIN vccd_1p0.gds1027
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 23.033 6.582 23.233 ;
 END
 END vccd_1p0.gds1027
 PIN vccd_1p0.gds1028
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.6 24.322 5.656 24.522 ;
 RECT 5.432 24.2335 5.488 24.4335 ;
 RECT 5.264 24.322 5.32 24.522 ;
 RECT 5.936 24.2335 5.992 24.4335 ;
 RECT 5.768 24.2335 5.824 24.4335 ;
 RECT 6.44 24.2505 6.496 24.4505 ;
 RECT 6.272 24.2335 6.328 24.4335 ;
 RECT 6.104 24.322 6.16 24.522 ;
 RECT 5.6 23.062 5.656 23.262 ;
 RECT 5.432 22.9735 5.488 23.1735 ;
 RECT 5.264 23.062 5.32 23.262 ;
 RECT 5.936 22.9735 5.992 23.1735 ;
 RECT 5.768 22.9735 5.824 23.1735 ;
 RECT 6.44 22.9905 6.496 23.1905 ;
 RECT 6.272 22.9735 6.328 23.1735 ;
 RECT 6.104 23.062 6.16 23.262 ;
 RECT 5.6 21.802 5.656 22.002 ;
 RECT 5.432 21.7135 5.488 21.9135 ;
 RECT 5.264 21.802 5.32 22.002 ;
 RECT 5.936 21.7135 5.992 21.9135 ;
 RECT 5.768 21.7135 5.824 21.9135 ;
 RECT 6.44 21.7305 6.496 21.9305 ;
 RECT 6.272 21.7135 6.328 21.9135 ;
 RECT 6.104 21.802 6.16 22.002 ;
 RECT 5.6 20.542 5.656 20.742 ;
 RECT 5.264 20.542 5.32 20.742 ;
 RECT 5.432 20.4535 5.488 20.6535 ;
 RECT 5.768 20.4535 5.824 20.6535 ;
 RECT 5.936 20.4535 5.992 20.6535 ;
 RECT 6.44 20.4705 6.496 20.6705 ;
 RECT 6.104 20.542 6.16 20.742 ;
 RECT 6.272 20.4535 6.328 20.6535 ;
 END
 END vccd_1p0.gds1028
 PIN vccd_1p0.gds1029
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 20.764 13.978 20.964 ;
 END
 END vccd_1p0.gds1029
 PIN vccd_1p0.gds1030
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 23.284 13.978 23.484 ;
 END
 END vccd_1p0.gds1030
 PIN vccd_1p0.gds1031
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 22.024 13.978 22.224 ;
 END
 END vccd_1p0.gds1031
 PIN vccd_1p0.gds1032
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 24.544 13.978 24.744 ;
 END
 END vccd_1p0.gds1032
 PIN vccd_1p0.gds1033
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 24.544 14.398 24.744 ;
 END
 END vccd_1p0.gds1033
 PIN vccd_1p0.gds1034
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 24.6715 14.934 24.8715 ;
 END
 END vccd_1p0.gds1034
 PIN vccd_1p0.gds1035
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 22.024 14.398 22.224 ;
 END
 END vccd_1p0.gds1035
 PIN vccd_1p0.gds1036
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 22.1515 14.934 22.3515 ;
 END
 END vccd_1p0.gds1036
 PIN vccd_1p0.gds1037
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 23.284 14.398 23.484 ;
 END
 END vccd_1p0.gds1037
 PIN vccd_1p0.gds1038
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 23.4115 14.934 23.6115 ;
 END
 END vccd_1p0.gds1038
 PIN vccd_1p0.gds1039
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 20.764 14.398 20.964 ;
 END
 END vccd_1p0.gds1039
 PIN vccd_1p0.gds1040
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 20.8915 14.934 21.0915 ;
 END
 END vccd_1p0.gds1040
 PIN vccd_1p0.gds1041
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 23.904 13.738 24.104 ;
 END
 END vccd_1p0.gds1041
 PIN vccd_1p0.gds1042
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 24.1915 13.138 24.3915 ;
 END
 END vccd_1p0.gds1042
 PIN vccd_1p0.gds1043
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 22.676 12.898 22.876 ;
 END
 END vccd_1p0.gds1043
 PIN vccd_1p0.gds1044
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 21.846 14.742 22.046 ;
 END
 END vccd_1p0.gds1044
 PIN vccd_1p0.gds1045
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 23.47 12.654 23.67 ;
 END
 END vccd_1p0.gds1045
 PIN vccd_1p0.gds1046
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 20.9765 12.526 21.1765 ;
 END
 END vccd_1p0.gds1046
 PIN vccd_1p0.gds1047
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 20.828 16.226 21.028 ;
 END
 END vccd_1p0.gds1047
 PIN vccd_1p0.gds1048
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 23.348 16.226 23.548 ;
 END
 END vccd_1p0.gds1048
 PIN vccd_1p0.gds1049
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 24.608 16.226 24.808 ;
 END
 END vccd_1p0.gds1049
 PIN vccd_1p0.gds1050
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 22.088 16.226 22.288 ;
 END
 END vccd_1p0.gds1050
 PIN vccd_1p0.gds1051
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 23.718 15.742 23.918 ;
 END
 END vccd_1p0.gds1051
 PIN vccd_1p0.gds1052
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 24.786 15.29 24.986 ;
 END
 END vccd_1p0.gds1052
 PIN vccd_1p0.gds1053
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 24.6185 18.09 24.8185 ;
 END
 END vccd_1p0.gds1053
 PIN vccd_1p0.gds1054
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 24.73 17.962 24.93 ;
 END
 END vccd_1p0.gds1054
 PIN vccd_1p0.gds1055
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 23.403 15.498 23.603 ;
 END
 END vccd_1p0.gds1055
 PIN vccd_1p0.gds1056
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 24.4565 17.734 24.6565 ;
 END
 END vccd_1p0.gds1056
 PIN vccd_1p0.gds1057
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 22.637 17.574 22.837 ;
 END
 END vccd_1p0.gds1057
 PIN vccd_1p0.gds1058
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 21.9335 17.154 22.1335 ;
 END
 END vccd_1p0.gds1058
 PIN vccd_1p0.gds1059
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 23.0125 23.842 23.2125 ;
 END
 END vccd_1p0.gds1059
 PIN vccd_1p0.gds1060
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 22.676 29.95 22.876 ;
 END
 END vccd_1p0.gds1060
 PIN vccd_1p0.gds1061
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 23.47 29.706 23.67 ;
 END
 END vccd_1p0.gds1061
 PIN vccd_1p0.gds1062
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 20.9765 29.578 21.1765 ;
 END
 END vccd_1p0.gds1062
 PIN vccd_1p0.gds1063
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 20.764 31.03 20.964 ;
 END
 END vccd_1p0.gds1063
 PIN vccd_1p0.gds1064
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 20.828 33.278 21.028 ;
 END
 END vccd_1p0.gds1064
 PIN vccd_1p0.gds1065
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 24.608 33.278 24.808 ;
 END
 END vccd_1p0.gds1065
 PIN vccd_1p0.gds1066
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 24.544 31.45 24.744 ;
 END
 END vccd_1p0.gds1066
 PIN vccd_1p0.gds1067
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 24.6715 31.986 24.8715 ;
 END
 END vccd_1p0.gds1067
 PIN vccd_1p0.gds1068
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 23.348 33.278 23.548 ;
 END
 END vccd_1p0.gds1068
 PIN vccd_1p0.gds1069
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 23.284 31.45 23.484 ;
 END
 END vccd_1p0.gds1069
 PIN vccd_1p0.gds1070
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 23.4115 31.986 23.6115 ;
 END
 END vccd_1p0.gds1070
 PIN vccd_1p0.gds1071
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 22.088 33.278 22.288 ;
 END
 END vccd_1p0.gds1071
 PIN vccd_1p0.gds1072
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 22.024 31.45 22.224 ;
 END
 END vccd_1p0.gds1072
 PIN vccd_1p0.gds1073
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 22.1515 31.986 22.3515 ;
 END
 END vccd_1p0.gds1073
 PIN vccd_1p0.gds1074
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 23.718 32.794 23.918 ;
 END
 END vccd_1p0.gds1074
 PIN vccd_1p0.gds1075
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 24.786 32.342 24.986 ;
 END
 END vccd_1p0.gds1075
 PIN vccd_1p0.gds1076
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 20.764 31.45 20.964 ;
 END
 END vccd_1p0.gds1076
 PIN vccd_1p0.gds1077
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 20.8915 31.986 21.0915 ;
 END
 END vccd_1p0.gds1077
 PIN vccd_1p0.gds1078
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 23.284 31.03 23.484 ;
 END
 END vccd_1p0.gds1078
 PIN vccd_1p0.gds1079
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 22.024 31.03 22.224 ;
 END
 END vccd_1p0.gds1079
 PIN vccd_1p0.gds1080
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 23.904 30.79 24.104 ;
 END
 END vccd_1p0.gds1080
 PIN vccd_1p0.gds1081
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 24.544 31.03 24.744 ;
 END
 END vccd_1p0.gds1081
 PIN vccd_1p0.gds1082
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 24.1915 30.19 24.3915 ;
 END
 END vccd_1p0.gds1082
 PIN vccd_1p0.gds1083
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 21.846 31.794 22.046 ;
 END
 END vccd_1p0.gds1083
 PIN vccd_1p0.gds1084
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 24.6185 35.142 24.8185 ;
 END
 END vccd_1p0.gds1084
 PIN vccd_1p0.gds1085
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 24.73 35.014 24.93 ;
 END
 END vccd_1p0.gds1085
 PIN vccd_1p0.gds1086
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 23.403 32.55 23.603 ;
 END
 END vccd_1p0.gds1086
 PIN vccd_1p0.gds1087
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 24.44 34.786 24.64 ;
 END
 END vccd_1p0.gds1087
 PIN vccd_1p0.gds1088
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 22.6315 34.626 22.8315 ;
 END
 END vccd_1p0.gds1088
 PIN vccd_1p0.gds1089
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 21.9335 34.206 22.1335 ;
 END
 END vccd_1p0.gds1089
 PIN vccd_1p0.gds1090
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 23.0125 40.894 23.2125 ;
 END
 END vccd_1p0.gds1090
 PIN vccd_1p0.gds1091
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 20.764 48.082 20.964 ;
 END
 END vccd_1p0.gds1091
 PIN vccd_1p0.gds1092
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 22.024 48.082 22.224 ;
 END
 END vccd_1p0.gds1092
 PIN vccd_1p0.gds1093
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 24.544 48.502 24.744 ;
 END
 END vccd_1p0.gds1093
 PIN vccd_1p0.gds1094
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 24.6715 49.038 24.8715 ;
 END
 END vccd_1p0.gds1094
 PIN vccd_1p0.gds1095
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 23.284 48.502 23.484 ;
 END
 END vccd_1p0.gds1095
 PIN vccd_1p0.gds1096
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 23.4115 49.038 23.6115 ;
 END
 END vccd_1p0.gds1096
 PIN vccd_1p0.gds1097
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 22.024 48.502 22.224 ;
 END
 END vccd_1p0.gds1097
 PIN vccd_1p0.gds1098
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 22.1515 49.038 22.3515 ;
 END
 END vccd_1p0.gds1098
 PIN vccd_1p0.gds1099
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 23.718 49.846 23.918 ;
 END
 END vccd_1p0.gds1099
 PIN vccd_1p0.gds1100
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 24.786 49.394 24.986 ;
 END
 END vccd_1p0.gds1100
 PIN vccd_1p0.gds1101
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 20.764 48.502 20.964 ;
 END
 END vccd_1p0.gds1101
 PIN vccd_1p0.gds1102
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 20.8915 49.038 21.0915 ;
 END
 END vccd_1p0.gds1102
 PIN vccd_1p0.gds1103
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 24.544 48.082 24.744 ;
 END
 END vccd_1p0.gds1103
 PIN vccd_1p0.gds1104
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 23.904 47.842 24.104 ;
 END
 END vccd_1p0.gds1104
 PIN vccd_1p0.gds1105
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 23.284 48.082 23.484 ;
 END
 END vccd_1p0.gds1105
 PIN vccd_1p0.gds1106
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 24.1915 47.242 24.3915 ;
 END
 END vccd_1p0.gds1106
 PIN vccd_1p0.gds1107
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 22.676 47.002 22.876 ;
 END
 END vccd_1p0.gds1107
 PIN vccd_1p0.gds1108
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 21.846 48.846 22.046 ;
 END
 END vccd_1p0.gds1108
 PIN vccd_1p0.gds1109
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 23.403 49.602 23.603 ;
 END
 END vccd_1p0.gds1109
 PIN vccd_1p0.gds1110
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 23.47 46.758 23.67 ;
 END
 END vccd_1p0.gds1110
 PIN vccd_1p0.gds1111
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 20.9765 46.63 21.1765 ;
 END
 END vccd_1p0.gds1111
 PIN vccd_1p0.gds1112
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 20.828 50.33 21.028 ;
 END
 END vccd_1p0.gds1112
 PIN vccd_1p0.gds1113
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 24.608 50.33 24.808 ;
 END
 END vccd_1p0.gds1113
 PIN vccd_1p0.gds1114
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 23.348 50.33 23.548 ;
 END
 END vccd_1p0.gds1114
 PIN vccd_1p0.gds1115
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 22.088 50.33 22.288 ;
 END
 END vccd_1p0.gds1115
 PIN vccd_1p0.gds1116
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 22.637 51.678 22.837 ;
 END
 END vccd_1p0.gds1116
 PIN vccd_1p0.gds1117
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 24.6185 52.194 24.8185 ;
 END
 END vccd_1p0.gds1117
 PIN vccd_1p0.gds1118
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 24.73 52.066 24.93 ;
 END
 END vccd_1p0.gds1118
 PIN vccd_1p0.gds1119
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 21.9335 51.258 22.1335 ;
 END
 END vccd_1p0.gds1119
 PIN vccd_1p0.gds1120
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 24.4565 51.838 24.6565 ;
 END
 END vccd_1p0.gds1120
 PIN vccd_1p0.gds1121
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 23.0125 57.946 23.2125 ;
 END
 END vccd_1p0.gds1121
 PIN vccd_1p0.gds1122
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 20.764 65.134 20.964 ;
 END
 END vccd_1p0.gds1122
 PIN vccd_1p0.gds1123
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 22.024 65.134 22.224 ;
 END
 END vccd_1p0.gds1123
 PIN vccd_1p0.gds1124
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 24.544 65.134 24.744 ;
 END
 END vccd_1p0.gds1124
 PIN vccd_1p0.gds1125
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 23.904 64.894 24.104 ;
 END
 END vccd_1p0.gds1125
 PIN vccd_1p0.gds1126
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 23.284 65.134 23.484 ;
 END
 END vccd_1p0.gds1126
 PIN vccd_1p0.gds1127
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 24.1915 64.294 24.3915 ;
 END
 END vccd_1p0.gds1127
 PIN vccd_1p0.gds1128
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 23.47 63.81 23.67 ;
 END
 END vccd_1p0.gds1128
 PIN vccd_1p0.gds1129
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 20.9765 63.682 21.1765 ;
 END
 END vccd_1p0.gds1129
 PIN vccd_1p0.gds1130
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 22.676 64.054 22.876 ;
 END
 END vccd_1p0.gds1130
 PIN vccd_1p0.gds1131
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 20.828 67.382 21.028 ;
 END
 END vccd_1p0.gds1131
 PIN vccd_1p0.gds1132
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 22.088 67.382 22.288 ;
 END
 END vccd_1p0.gds1132
 PIN vccd_1p0.gds1133
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 22.024 65.554 22.224 ;
 END
 END vccd_1p0.gds1133
 PIN vccd_1p0.gds1134
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 22.1515 66.09 22.3515 ;
 END
 END vccd_1p0.gds1134
 PIN vccd_1p0.gds1135
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 23.348 67.382 23.548 ;
 END
 END vccd_1p0.gds1135
 PIN vccd_1p0.gds1136
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 23.284 65.554 23.484 ;
 END
 END vccd_1p0.gds1136
 PIN vccd_1p0.gds1137
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 23.4115 66.09 23.6115 ;
 END
 END vccd_1p0.gds1137
 PIN vccd_1p0.gds1138
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 24.608 67.382 24.808 ;
 END
 END vccd_1p0.gds1138
 PIN vccd_1p0.gds1139
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 24.544 65.554 24.744 ;
 END
 END vccd_1p0.gds1139
 PIN vccd_1p0.gds1140
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 24.6715 66.09 24.8715 ;
 END
 END vccd_1p0.gds1140
 PIN vccd_1p0.gds1141
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 24.786 66.446 24.986 ;
 END
 END vccd_1p0.gds1141
 PIN vccd_1p0.gds1142
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 20.764 65.554 20.964 ;
 END
 END vccd_1p0.gds1142
 PIN vccd_1p0.gds1143
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 20.8915 66.09 21.0915 ;
 END
 END vccd_1p0.gds1143
 PIN vccd_1p0.gds1144
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 21.846 65.898 22.046 ;
 END
 END vccd_1p0.gds1144
 PIN vccd_1p0.gds1145
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 22.637 68.73 22.837 ;
 END
 END vccd_1p0.gds1145
 PIN vccd_1p0.gds1146
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 24.6185 69.246 24.8185 ;
 END
 END vccd_1p0.gds1146
 PIN vccd_1p0.gds1147
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 24.73 69.118 24.93 ;
 END
 END vccd_1p0.gds1147
 PIN vccd_1p0.gds1148
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 21.9335 68.31 22.1335 ;
 END
 END vccd_1p0.gds1148
 PIN vccd_1p0.gds1149
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 23.403 66.654 23.603 ;
 END
 END vccd_1p0.gds1149
 PIN vccd_1p0.gds1150
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 24.4565 68.89 24.6565 ;
 END
 END vccd_1p0.gds1150
 PIN vccd_1p0.gds1151
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 23.718 66.898 23.918 ;
 END
 END vccd_1p0.gds1151
 PIN vccd_1p0.gds1152
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 27.163 0.43 27.363 ;
 END
 END vccd_1p0.gds1152
 PIN vccd_1p0.gds1153
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 27.949 5.202 28.149 ;
 END
 END vccd_1p0.gds1153
 PIN vccd_1p0.gds1154
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 27.977 1.542 28.177 ;
 END
 END vccd_1p0.gds1154
 PIN vccd_1p0.gds1155
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 26.717 1.542 26.917 ;
 END
 END vccd_1p0.gds1155
 PIN vccd_1p0.gds1156
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 27.3585 0.548 27.5585 ;
 END
 END vccd_1p0.gds1156
 PIN vccd_1p0.gds1157
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 25.457 1.542 25.657 ;
 END
 END vccd_1p0.gds1157
 PIN vccd_1p0.gds1158
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 27.1755 0.858 27.3755 ;
 END
 END vccd_1p0.gds1158
 PIN vccd_1p0.gds1159
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 27.154 1.362 27.354 ;
 END
 END vccd_1p0.gds1159
 PIN vccd_1p0.gds1160
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 27.1375 1.218 27.3375 ;
 END
 END vccd_1p0.gds1160
 PIN vccd_1p0.gds1161
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 27.166 1.09 27.366 ;
 END
 END vccd_1p0.gds1161
 PIN vccd_1p0.gds1162
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 27.9065 1.782 28.1065 ;
 END
 END vccd_1p0.gds1162
 PIN vccd_1p0.gds1163
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 28.168 2.202 28.368 ;
 END
 END vccd_1p0.gds1163
 PIN vccd_1p0.gds1164
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 27.051 2.622 27.251 ;
 END
 END vccd_1p0.gds1164
 PIN vccd_1p0.gds1165
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 26.5995 5.202 26.7995 ;
 END
 END vccd_1p0.gds1165
 PIN vccd_1p0.gds1166
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 28.5475 3.666 28.7475 ;
 END
 END vccd_1p0.gds1166
 PIN vccd_1p0.gds1167
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 25.9265 3.666 26.1265 ;
 END
 END vccd_1p0.gds1167
 PIN vccd_1p0.gds1168
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 28.527 4.738 28.727 ;
 END
 END vccd_1p0.gds1168
 PIN vccd_1p0.gds1169
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 25.9915 4.738 26.1915 ;
 END
 END vccd_1p0.gds1169
 PIN vccd_1p0.gds1170
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 28.2865 2.462 28.4865 ;
 END
 END vccd_1p0.gds1170
 PIN vccd_1p0.gds1171
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 26.9365 1.962 27.1365 ;
 END
 END vccd_1p0.gds1171
 PIN vccd_1p0.gds1172
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 27.0225 3.042 27.2225 ;
 END
 END vccd_1p0.gds1172
 PIN vccd_1p0.gds1173
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 27.098 2.882 27.298 ;
 END
 END vccd_1p0.gds1173
 PIN vccd_1p0.gds1174
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 27.1435 3.262 27.3435 ;
 END
 END vccd_1p0.gds1174
 PIN vccd_1p0.gds1175
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 27.1225 3.39 27.3225 ;
 END
 END vccd_1p0.gds1175
 PIN vccd_1p0.gds1176
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 27.157 3.858 27.357 ;
 END
 END vccd_1p0.gds1176
 PIN vccd_1p0.gds1177
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 26.4645 4.258 26.6645 ;
 END
 END vccd_1p0.gds1177
 PIN vccd_1p0.gds1178
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 28.42 4.066 28.62 ;
 END
 END vccd_1p0.gds1178
 PIN vccd_1p0.gds1179
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 25.5365 4.066 25.7365 ;
 END
 END vccd_1p0.gds1179
 PIN vccd_1p0.gds1180
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 27.148 4.546 27.348 ;
 END
 END vccd_1p0.gds1180
 PIN vccd_1p0.gds1181
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 27.1645 5.01 27.3645 ;
 END
 END vccd_1p0.gds1181
 PIN vccd_1p0.gds1182
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 3.584 28.0035 3.64 28.2035 ;
 RECT 3.584 26.7435 3.64 26.9435 ;
 RECT 3.584 25.4835 3.64 25.6835 ;
 RECT 4.34 28.102 4.396 28.302 ;
 RECT 4.172 28.102 4.228 28.302 ;
 RECT 4.76 28.0615 4.816 28.2615 ;
 RECT 5.096 28.102 5.152 28.302 ;
 RECT 4.928 28.0615 4.984 28.2615 ;
 RECT 4.34 26.842 4.396 27.042 ;
 RECT 4.172 26.842 4.228 27.042 ;
 RECT 4.76 26.8015 4.816 27.0015 ;
 RECT 5.096 26.842 5.152 27.042 ;
 RECT 4.928 26.8015 4.984 27.0015 ;
 RECT 4.34 25.582 4.396 25.782 ;
 RECT 4.172 25.582 4.228 25.782 ;
 RECT 4.76 25.5415 4.816 25.7415 ;
 RECT 5.096 25.582 5.152 25.782 ;
 RECT 4.928 25.5415 4.984 25.7415 ;
 END
 END vccd_1p0.gds1182
 PIN vccd_1p0.gds1183
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 27.157 6.838 27.357 ;
 END
 END vccd_1p0.gds1183
 PIN vccd_1p0.gds1184
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 28.3495 6.05 28.5495 ;
 END
 END vccd_1p0.gds1184
 PIN vccd_1p0.gds1185
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.754 26.2565 5.794 26.4565 ;
 END
 END vccd_1p0.gds1185
 PIN vccd_1p0.gds1186
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 28.5475 5.41 28.7475 ;
 END
 END vccd_1p0.gds1186
 PIN vccd_1p0.gds1187
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 25.8965 5.41 26.0965 ;
 END
 END vccd_1p0.gds1187
 PIN vccd_1p0.gds1188
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 28.094 5.922 28.294 ;
 END
 END vccd_1p0.gds1188
 PIN vccd_1p0.gds1189
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 27.165 5.602 27.365 ;
 END
 END vccd_1p0.gds1189
 PIN vccd_1p0.gds1190
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 27.696 6.306 27.896 ;
 END
 END vccd_1p0.gds1190
 PIN vccd_1p0.gds1191
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 27.129 6.582 27.329 ;
 END
 END vccd_1p0.gds1191
 PIN vccd_1p0.gds1192
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.6 28.102 5.656 28.302 ;
 RECT 5.432 28.0135 5.488 28.2135 ;
 RECT 5.264 28.102 5.32 28.302 ;
 RECT 5.936 28.0135 5.992 28.2135 ;
 RECT 5.768 28.0135 5.824 28.2135 ;
 RECT 6.44 28.0305 6.496 28.2305 ;
 RECT 6.272 28.0135 6.328 28.2135 ;
 RECT 6.104 28.102 6.16 28.302 ;
 RECT 5.6 26.842 5.656 27.042 ;
 RECT 5.432 26.7535 5.488 26.9535 ;
 RECT 5.264 26.842 5.32 27.042 ;
 RECT 5.936 26.7535 5.992 26.9535 ;
 RECT 5.768 26.7535 5.824 26.9535 ;
 RECT 6.44 26.7705 6.496 26.9705 ;
 RECT 6.272 26.7535 6.328 26.9535 ;
 RECT 6.104 26.842 6.16 27.042 ;
 RECT 5.6 25.582 5.656 25.782 ;
 RECT 5.432 25.4935 5.488 25.6935 ;
 RECT 5.264 25.582 5.32 25.782 ;
 RECT 5.936 25.4935 5.992 25.6935 ;
 RECT 5.768 25.4935 5.824 25.6935 ;
 RECT 6.44 25.5105 6.496 25.7105 ;
 RECT 6.272 25.4935 6.328 25.6935 ;
 RECT 6.104 25.582 6.16 25.782 ;
 END
 END vccd_1p0.gds1192
 PIN vccd_1p0.gds1193
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 27.064 13.978 27.264 ;
 END
 END vccd_1p0.gds1193
 PIN vccd_1p0.gds1194
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 28.324 13.978 28.524 ;
 END
 END vccd_1p0.gds1194
 PIN vccd_1p0.gds1195
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 25.804 13.978 26.004 ;
 END
 END vccd_1p0.gds1195
 PIN vccd_1p0.gds1196
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 27.064 14.398 27.264 ;
 END
 END vccd_1p0.gds1196
 PIN vccd_1p0.gds1197
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 25.804 14.398 26.004 ;
 END
 END vccd_1p0.gds1197
 PIN vccd_1p0.gds1198
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 25.9315 14.934 26.1315 ;
 END
 END vccd_1p0.gds1198
 PIN vccd_1p0.gds1199
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 28.324 14.398 28.524 ;
 END
 END vccd_1p0.gds1199
 PIN vccd_1p0.gds1200
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 28.4515 14.934 28.6515 ;
 END
 END vccd_1p0.gds1200
 PIN vccd_1p0.gds1201
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 27.454 13.738 27.654 ;
 END
 END vccd_1p0.gds1201
 PIN vccd_1p0.gds1202
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 27.6475 13.138 27.8475 ;
 END
 END vccd_1p0.gds1202
 PIN vccd_1p0.gds1203
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 26.9635 12.898 27.1635 ;
 END
 END vccd_1p0.gds1203
 PIN vccd_1p0.gds1204
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 26.562 14.742 26.762 ;
 END
 END vccd_1p0.gds1204
 PIN vccd_1p0.gds1205
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 27.1915 14.934 27.3915 ;
 END
 END vccd_1p0.gds1205
 PIN vccd_1p0.gds1206
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 27.3545 12.654 27.5545 ;
 END
 END vccd_1p0.gds1206
 PIN vccd_1p0.gds1207
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 28.5475 12.526 28.7475 ;
 END
 END vccd_1p0.gds1207
 PIN vccd_1p0.gds1208
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 25.948 12.526 26.148 ;
 END
 END vccd_1p0.gds1208
 PIN vccd_1p0.gds1209
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 27.128 16.226 27.328 ;
 END
 END vccd_1p0.gds1209
 PIN vccd_1p0.gds1210
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 28.388 16.226 28.588 ;
 END
 END vccd_1p0.gds1210
 PIN vccd_1p0.gds1211
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 25.868 16.226 26.068 ;
 END
 END vccd_1p0.gds1211
 PIN vccd_1p0.gds1212
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 27.498 15.742 27.698 ;
 END
 END vccd_1p0.gds1212
 PIN vccd_1p0.gds1213
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 28.032 15.29 28.232 ;
 END
 END vccd_1p0.gds1213
 PIN vccd_1p0.gds1214
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 27.91 18.09 28.11 ;
 END
 END vccd_1p0.gds1214
 PIN vccd_1p0.gds1215
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 27.984 17.962 28.184 ;
 END
 END vccd_1p0.gds1215
 PIN vccd_1p0.gds1216
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 27.3415 15.498 27.5415 ;
 END
 END vccd_1p0.gds1216
 PIN vccd_1p0.gds1217
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 27.8695 17.734 28.0695 ;
 END
 END vccd_1p0.gds1217
 PIN vccd_1p0.gds1218
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 26.904 17.574 27.104 ;
 END
 END vccd_1p0.gds1218
 PIN vccd_1p0.gds1219
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 26.5335 17.154 26.7335 ;
 END
 END vccd_1p0.gds1219
 PIN vccd_1p0.gds1220
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 27.1095 23.842 27.3095 ;
 END
 END vccd_1p0.gds1220
 PIN vccd_1p0.gds1221
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 26.9635 29.95 27.1635 ;
 END
 END vccd_1p0.gds1221
 PIN vccd_1p0.gds1222
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 27.3545 29.706 27.5545 ;
 END
 END vccd_1p0.gds1222
 PIN vccd_1p0.gds1223
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 28.5475 29.578 28.7475 ;
 END
 END vccd_1p0.gds1223
 PIN vccd_1p0.gds1224
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 25.948 29.578 26.148 ;
 END
 END vccd_1p0.gds1224
 PIN vccd_1p0.gds1225
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 27.064 31.03 27.264 ;
 END
 END vccd_1p0.gds1225
 PIN vccd_1p0.gds1226
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 27.128 33.278 27.328 ;
 END
 END vccd_1p0.gds1226
 PIN vccd_1p0.gds1227
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 27.064 31.45 27.264 ;
 END
 END vccd_1p0.gds1227
 PIN vccd_1p0.gds1228
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 28.388 33.278 28.588 ;
 END
 END vccd_1p0.gds1228
 PIN vccd_1p0.gds1229
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 25.868 33.278 26.068 ;
 END
 END vccd_1p0.gds1229
 PIN vccd_1p0.gds1230
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 27.498 32.794 27.698 ;
 END
 END vccd_1p0.gds1230
 PIN vccd_1p0.gds1231
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 25.804 31.45 26.004 ;
 END
 END vccd_1p0.gds1231
 PIN vccd_1p0.gds1232
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 25.9315 31.986 26.1315 ;
 END
 END vccd_1p0.gds1232
 PIN vccd_1p0.gds1233
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 28.032 32.342 28.232 ;
 END
 END vccd_1p0.gds1233
 PIN vccd_1p0.gds1234
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 28.324 31.03 28.524 ;
 END
 END vccd_1p0.gds1234
 PIN vccd_1p0.gds1235
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 25.804 31.03 26.004 ;
 END
 END vccd_1p0.gds1235
 PIN vccd_1p0.gds1236
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 27.454 30.79 27.654 ;
 END
 END vccd_1p0.gds1236
 PIN vccd_1p0.gds1237
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 27.6475 30.19 27.8475 ;
 END
 END vccd_1p0.gds1237
 PIN vccd_1p0.gds1238
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 26.562 31.794 26.762 ;
 END
 END vccd_1p0.gds1238
 PIN vccd_1p0.gds1239
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 28.324 31.45 28.524 ;
 END
 END vccd_1p0.gds1239
 PIN vccd_1p0.gds1240
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 28.4515 31.986 28.6515 ;
 END
 END vccd_1p0.gds1240
 PIN vccd_1p0.gds1241
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 27.91 35.142 28.11 ;
 END
 END vccd_1p0.gds1241
 PIN vccd_1p0.gds1242
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 27.984 35.014 28.184 ;
 END
 END vccd_1p0.gds1242
 PIN vccd_1p0.gds1243
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 27.1915 31.986 27.3915 ;
 END
 END vccd_1p0.gds1243
 PIN vccd_1p0.gds1244
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 27.3415 32.55 27.5415 ;
 END
 END vccd_1p0.gds1244
 PIN vccd_1p0.gds1245
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 27.845 34.786 28.045 ;
 END
 END vccd_1p0.gds1245
 PIN vccd_1p0.gds1246
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 26.926 34.626 27.126 ;
 END
 END vccd_1p0.gds1246
 PIN vccd_1p0.gds1247
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 26.5335 34.206 26.7335 ;
 END
 END vccd_1p0.gds1247
 PIN vccd_1p0.gds1248
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 27.1095 40.894 27.3095 ;
 END
 END vccd_1p0.gds1248
 PIN vccd_1p0.gds1249
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 27.064 48.082 27.264 ;
 END
 END vccd_1p0.gds1249
 PIN vccd_1p0.gds1250
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 28.324 48.082 28.524 ;
 END
 END vccd_1p0.gds1250
 PIN vccd_1p0.gds1251
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 25.804 48.082 26.004 ;
 END
 END vccd_1p0.gds1251
 PIN vccd_1p0.gds1252
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 27.064 48.502 27.264 ;
 END
 END vccd_1p0.gds1252
 PIN vccd_1p0.gds1253
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 27.498 49.846 27.698 ;
 END
 END vccd_1p0.gds1253
 PIN vccd_1p0.gds1254
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 25.804 48.502 26.004 ;
 END
 END vccd_1p0.gds1254
 PIN vccd_1p0.gds1255
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 25.9315 49.038 26.1315 ;
 END
 END vccd_1p0.gds1255
 PIN vccd_1p0.gds1256
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 28.032 49.394 28.232 ;
 END
 END vccd_1p0.gds1256
 PIN vccd_1p0.gds1257
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 27.454 47.842 27.654 ;
 END
 END vccd_1p0.gds1257
 PIN vccd_1p0.gds1258
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 27.6475 47.242 27.8475 ;
 END
 END vccd_1p0.gds1258
 PIN vccd_1p0.gds1259
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 26.9635 47.002 27.1635 ;
 END
 END vccd_1p0.gds1259
 PIN vccd_1p0.gds1260
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 26.562 48.846 26.762 ;
 END
 END vccd_1p0.gds1260
 PIN vccd_1p0.gds1261
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 28.324 48.502 28.524 ;
 END
 END vccd_1p0.gds1261
 PIN vccd_1p0.gds1262
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 28.4515 49.038 28.6515 ;
 END
 END vccd_1p0.gds1262
 PIN vccd_1p0.gds1263
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 27.1915 49.038 27.3915 ;
 END
 END vccd_1p0.gds1263
 PIN vccd_1p0.gds1264
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 27.3415 49.602 27.5415 ;
 END
 END vccd_1p0.gds1264
 PIN vccd_1p0.gds1265
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 27.3545 46.758 27.5545 ;
 END
 END vccd_1p0.gds1265
 PIN vccd_1p0.gds1266
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 28.5475 46.63 28.7475 ;
 END
 END vccd_1p0.gds1266
 PIN vccd_1p0.gds1267
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 25.948 46.63 26.148 ;
 END
 END vccd_1p0.gds1267
 PIN vccd_1p0.gds1268
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 27.128 50.33 27.328 ;
 END
 END vccd_1p0.gds1268
 PIN vccd_1p0.gds1269
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 28.388 50.33 28.588 ;
 END
 END vccd_1p0.gds1269
 PIN vccd_1p0.gds1270
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 25.868 50.33 26.068 ;
 END
 END vccd_1p0.gds1270
 PIN vccd_1p0.gds1271
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 26.904 51.678 27.104 ;
 END
 END vccd_1p0.gds1271
 PIN vccd_1p0.gds1272
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 27.91 52.194 28.11 ;
 END
 END vccd_1p0.gds1272
 PIN vccd_1p0.gds1273
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 27.984 52.066 28.184 ;
 END
 END vccd_1p0.gds1273
 PIN vccd_1p0.gds1274
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 26.5335 51.258 26.7335 ;
 END
 END vccd_1p0.gds1274
 PIN vccd_1p0.gds1275
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 27.8695 51.838 28.0695 ;
 END
 END vccd_1p0.gds1275
 PIN vccd_1p0.gds1276
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 27.1095 57.946 27.3095 ;
 END
 END vccd_1p0.gds1276
 PIN vccd_1p0.gds1277
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 27.064 65.134 27.264 ;
 END
 END vccd_1p0.gds1277
 PIN vccd_1p0.gds1278
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 28.324 65.134 28.524 ;
 END
 END vccd_1p0.gds1278
 PIN vccd_1p0.gds1279
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 25.804 65.134 26.004 ;
 END
 END vccd_1p0.gds1279
 PIN vccd_1p0.gds1280
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 27.454 64.894 27.654 ;
 END
 END vccd_1p0.gds1280
 PIN vccd_1p0.gds1281
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 27.6475 64.294 27.8475 ;
 END
 END vccd_1p0.gds1281
 PIN vccd_1p0.gds1282
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 27.3545 63.81 27.5545 ;
 END
 END vccd_1p0.gds1282
 PIN vccd_1p0.gds1283
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 28.5475 63.682 28.7475 ;
 END
 END vccd_1p0.gds1283
 PIN vccd_1p0.gds1284
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 25.948 63.682 26.148 ;
 END
 END vccd_1p0.gds1284
 PIN vccd_1p0.gds1285
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 26.9635 64.054 27.1635 ;
 END
 END vccd_1p0.gds1285
 PIN vccd_1p0.gds1286
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 27.128 67.382 27.328 ;
 END
 END vccd_1p0.gds1286
 PIN vccd_1p0.gds1287
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 27.064 65.554 27.264 ;
 END
 END vccd_1p0.gds1287
 PIN vccd_1p0.gds1288
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 28.388 67.382 28.588 ;
 END
 END vccd_1p0.gds1288
 PIN vccd_1p0.gds1289
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 25.868 67.382 26.068 ;
 END
 END vccd_1p0.gds1289
 PIN vccd_1p0.gds1290
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 25.804 65.554 26.004 ;
 END
 END vccd_1p0.gds1290
 PIN vccd_1p0.gds1291
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 25.9315 66.09 26.1315 ;
 END
 END vccd_1p0.gds1291
 PIN vccd_1p0.gds1292
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 28.032 66.446 28.232 ;
 END
 END vccd_1p0.gds1292
 PIN vccd_1p0.gds1293
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 26.562 65.898 26.762 ;
 END
 END vccd_1p0.gds1293
 PIN vccd_1p0.gds1294
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 28.324 65.554 28.524 ;
 END
 END vccd_1p0.gds1294
 PIN vccd_1p0.gds1295
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 28.4515 66.09 28.6515 ;
 END
 END vccd_1p0.gds1295
 PIN vccd_1p0.gds1296
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 26.904 68.73 27.104 ;
 END
 END vccd_1p0.gds1296
 PIN vccd_1p0.gds1297
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 27.91 69.246 28.11 ;
 END
 END vccd_1p0.gds1297
 PIN vccd_1p0.gds1298
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 27.984 69.118 28.184 ;
 END
 END vccd_1p0.gds1298
 PIN vccd_1p0.gds1299
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 26.5335 68.31 26.7335 ;
 END
 END vccd_1p0.gds1299
 PIN vccd_1p0.gds1300
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 27.1915 66.09 27.3915 ;
 END
 END vccd_1p0.gds1300
 PIN vccd_1p0.gds1301
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 27.3415 66.654 27.5415 ;
 END
 END vccd_1p0.gds1301
 PIN vccd_1p0.gds1302
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 27.8695 68.89 28.0695 ;
 END
 END vccd_1p0.gds1302
 PIN vccd_1p0.gds1303
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 27.498 66.898 27.698 ;
 END
 END vccd_1p0.gds1303
 PIN vss
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 0.913 2.962 1.113 ;
 END
 END vss
 PIN vss.gds1
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 2.294 0.29 2.494 ;
 END
 END vss.gds1
 PIN vss.gds2
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 2.173 2.962 2.373 ;
 END
 END vss.gds2
 PIN vss.gds3
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 3.433 2.962 3.633 ;
 END
 END vss.gds3
 PIN vss.gds4
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 4.693 2.962 4.893 ;
 END
 END vss.gds4
 PIN vss.gds5
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 0.6075 3.142 0.8075 ;
 END
 END vss.gds5
 PIN vss.gds6
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 4.292 3.142 4.492 ;
 END
 END vss.gds6
 PIN vss.gds7
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.286 2.803 3.326 3.003 ;
 END
 END vss.gds7
 PIN vss.gds8
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.754 2.803 3.794 3.003 ;
 END
 END vss.gds8
 PIN vss.gds9
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.442 2.397 4.482 2.597 ;
 END
 END vss.gds9
 PIN vss.gds10
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 2.598 0.602 2.798 ;
 END
 END vss.gds10
 PIN vss.gds11
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 1.772 3.142 1.972 ;
 END
 END vss.gds11
 PIN vss.gds12
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.414 3.079 3.454 3.279 ;
 END
 END vss.gds12
 PIN vss.gds13
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 2.397 0.942 2.597 ;
 END
 END vss.gds13
 PIN vss.gds14
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 2.941 1.282 3.141 ;
 END
 END vss.gds14
 PIN vss.gds15
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 2.8265 2.122 3.0265 ;
 END
 END vss.gds15
 PIN vss.gds16
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 2.397 4.882 2.597 ;
 END
 END vss.gds16
 PIN vss.gds17
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.57 2.6 4.61 2.8 ;
 END
 END vss.gds17
 PIN vss.gds18
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 2.803 4.194 3.003 ;
 END
 END vss.gds18
 PIN vss.gds19
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 2.803 5.074 3.003 ;
 END
 END vss.gds19
 PIN vss.gds20
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 3.032 3.142 3.232 ;
 END
 END vss.gds20
 PIN vss.gds21
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.562 3.079 3.602 3.279 ;
 END
 END vss.gds21
 PIN vss.gds22
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 2.6995 4.002 2.8995 ;
 END
 END vss.gds22
 PIN vss.gds23
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 2.6995 5.282 2.8995 ;
 END
 END vss.gds23
 PIN vss.gds24
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 2.738 2.302 2.938 ;
 END
 END vss.gds24
 PIN vss.gds25
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 3.1755 1.462 3.3755 ;
 END
 END vss.gds25
 PIN vss.gds26
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 2.4975 0.718 2.6975 ;
 END
 END vss.gds26
 PIN vss.gds27
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 2.576 0.9135 2.632 1.1135 ;
 RECT 2.408 0.9135 2.464 1.1135 ;
 RECT 2.996 0.9135 3.052 1.1135 ;
 RECT 3.332 1.005 3.388 1.205 ;
 RECT 3.5 0.9615 3.556 1.1615 ;
 RECT 0.98 0.8285 1.036 1.0285 ;
 RECT 2.072 0.829 2.128 1.029 ;
 RECT 2.576 2.1735 2.632 2.3735 ;
 RECT 2.408 2.1735 2.464 2.3735 ;
 RECT 2.996 2.1735 3.052 2.3735 ;
 RECT 3.332 2.265 3.388 2.465 ;
 RECT 3.5 2.2215 3.556 2.4215 ;
 RECT 0.98 2.0885 1.036 2.2885 ;
 RECT 2.072 2.089 2.128 2.289 ;
 RECT 2.576 3.4335 2.632 3.6335 ;
 RECT 2.408 3.4335 2.464 3.6335 ;
 RECT 2.996 3.4335 3.052 3.6335 ;
 RECT 3.332 3.525 3.388 3.725 ;
 RECT 3.5 3.4815 3.556 3.6815 ;
 RECT 0.98 3.3485 1.036 3.5485 ;
 RECT 2.072 3.349 2.128 3.549 ;
 RECT 2.576 4.6935 2.632 4.8935 ;
 RECT 2.408 4.6935 2.464 4.8935 ;
 RECT 2.996 4.6935 3.052 4.8935 ;
 RECT 3.332 4.785 3.388 4.985 ;
 RECT 3.5 4.7415 3.556 4.9415 ;
 RECT 0.98 4.6085 1.036 4.8085 ;
 RECT 2.072 4.609 2.128 4.809 ;
 RECT 0.392 4.699 0.448 4.899 ;
 RECT 0.812 4.785 0.868 4.985 ;
 RECT 0.644 4.699 0.7 4.899 ;
 RECT 1.232 4.699 1.288 4.899 ;
 RECT 1.4 4.699 1.456 4.899 ;
 RECT 1.568 4.699 1.624 4.899 ;
 RECT 1.82 4.699 1.876 4.899 ;
 RECT 2.24 4.699 2.296 4.899 ;
 RECT 2.744 4.609 2.8 4.809 ;
 RECT 3.164 4.699 3.22 4.899 ;
 RECT 3.92 4.699 3.976 4.899 ;
 RECT 3.752 4.969 3.808 5.169 ;
 RECT 4.508 4.8985 4.564 5.0985 ;
 RECT 0.392 3.439 0.448 3.639 ;
 RECT 0.812 3.525 0.868 3.725 ;
 RECT 0.644 3.439 0.7 3.639 ;
 RECT 1.232 3.439 1.288 3.639 ;
 RECT 1.4 3.439 1.456 3.639 ;
 RECT 1.568 3.439 1.624 3.639 ;
 RECT 1.82 3.439 1.876 3.639 ;
 RECT 2.24 3.439 2.296 3.639 ;
 RECT 2.744 3.349 2.8 3.549 ;
 RECT 3.164 3.439 3.22 3.639 ;
 RECT 3.92 3.439 3.976 3.639 ;
 RECT 3.752 3.709 3.808 3.909 ;
 RECT 4.508 3.6385 4.564 3.8385 ;
 RECT 0.392 2.179 0.448 2.379 ;
 RECT 0.812 2.265 0.868 2.465 ;
 RECT 0.644 2.179 0.7 2.379 ;
 RECT 1.232 2.179 1.288 2.379 ;
 RECT 1.4 2.179 1.456 2.379 ;
 RECT 1.568 2.179 1.624 2.379 ;
 RECT 1.82 2.179 1.876 2.379 ;
 RECT 2.24 2.179 2.296 2.379 ;
 RECT 2.744 2.089 2.8 2.289 ;
 RECT 3.164 2.179 3.22 2.379 ;
 RECT 3.92 2.179 3.976 2.379 ;
 RECT 3.752 2.449 3.808 2.649 ;
 RECT 4.508 2.3785 4.564 2.5785 ;
 RECT 0.392 0.919 0.448 1.119 ;
 RECT 0.812 1.005 0.868 1.205 ;
 RECT 0.644 0.919 0.7 1.119 ;
 RECT 1.232 0.919 1.288 1.119 ;
 RECT 1.4 0.919 1.456 1.119 ;
 RECT 1.568 0.919 1.624 1.119 ;
 RECT 1.82 0.919 1.876 1.119 ;
 RECT 2.24 0.919 2.296 1.119 ;
 RECT 2.744 0.829 2.8 1.029 ;
 RECT 3.164 0.919 3.22 1.119 ;
 RECT 3.92 0.919 3.976 1.119 ;
 RECT 3.752 1.189 3.808 1.389 ;
 RECT 4.508 1.1185 4.564 1.3185 ;
 END
 END vss.gds27
 PIN vss.gds28
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.134 3.0195 10.194 3.2195 ;
 END
 END vss.gds28
 PIN vss.gds29
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.966 3.0195 10.026 3.2195 ;
 END
 END vss.gds29
 PIN vss.gds30
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.798 3.0195 9.858 3.2195 ;
 END
 END vss.gds30
 PIN vss.gds31
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.79 3.0195 8.85 3.2195 ;
 END
 END vss.gds31
 PIN vss.gds32
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.622 3.0195 8.682 3.2195 ;
 END
 END vss.gds32
 PIN vss.gds33
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.454 3.0195 8.514 3.2195 ;
 END
 END vss.gds33
 PIN vss.gds34
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 3.0195 9.69 3.2195 ;
 END
 END vss.gds34
 PIN vss.gds35
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.118 3.0195 8.178 3.2195 ;
 END
 END vss.gds35
 PIN vss.gds36
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 3.0195 8.346 3.2195 ;
 END
 END vss.gds36
 PIN vss.gds37
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.95 3.0195 8.01 3.2195 ;
 END
 END vss.gds37
 PIN vss.gds38
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.782 3.0195 7.842 3.2195 ;
 END
 END vss.gds38
 PIN vss.gds39
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.462 3.0195 9.522 3.2195 ;
 END
 END vss.gds39
 PIN vss.gds40
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.294 3.0195 9.354 3.2195 ;
 END
 END vss.gds40
 PIN vss.gds41
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.126 3.0195 9.186 3.2195 ;
 END
 END vss.gds41
 PIN vss.gds42
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.446 3.0195 7.506 3.2195 ;
 END
 END vss.gds42
 PIN vss.gds43
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 3.0195 9.018 3.2195 ;
 END
 END vss.gds43
 PIN vss.gds44
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 3.0195 7.674 3.2195 ;
 END
 END vss.gds44
 PIN vss.gds45
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 2.803 5.474 3.003 ;
 END
 END vss.gds45
 PIN vss.gds46
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 2.803 5.986 3.003 ;
 END
 END vss.gds46
 PIN vss.gds47
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 2.803 5.73 3.003 ;
 END
 END vss.gds47
 PIN vss.gds48
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.278 3.0195 7.338 3.2195 ;
 END
 END vss.gds48
 PIN vss.gds49
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.11 3.0195 7.17 3.2195 ;
 END
 END vss.gds49
 PIN vss.gds50
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 2.599 6.434 2.799 ;
 END
 END vss.gds50
 PIN vss.gds51
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 2.6 6.178 2.8 ;
 END
 END vss.gds51
 PIN vss.gds52
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 6.524 4.661 6.58 4.861 ;
 RECT 6.524 3.401 6.58 3.601 ;
 RECT 6.524 2.141 6.58 2.341 ;
 RECT 6.692 4.984 6.748 5.184 ;
 RECT 6.692 3.724 6.748 3.924 ;
 RECT 6.692 2.464 6.748 2.664 ;
 RECT 6.692 1.204 6.748 1.404 ;
 RECT 6.608 4.969 6.664 5.169 ;
 RECT 6.608 3.709 6.664 3.909 ;
 RECT 6.608 2.449 6.664 2.649 ;
 RECT 6.608 1.189 6.664 1.389 ;
 RECT 6.524 0.881 6.58 1.081 ;
 END
 END vss.gds52
 PIN vss.gds53
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 1.458 14.87 1.658 ;
 END
 END vss.gds53
 PIN vss.gds54
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 2.678 13.898 2.878 ;
 END
 END vss.gds54
 PIN vss.gds55
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 2.718 14.87 2.918 ;
 END
 END vss.gds55
 PIN vss.gds56
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 3.938 13.898 4.138 ;
 END
 END vss.gds56
 PIN vss.gds57
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 3.978 14.87 4.178 ;
 END
 END vss.gds57
 PIN vss.gds58
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 5.198 13.898 5.398 ;
 END
 END vss.gds58
 PIN vss.gds59
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 5.238 14.87 5.438 ;
 END
 END vss.gds59
 PIN vss.gds60
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.15 3.0195 12.21 3.2195 ;
 END
 END vss.gds60
 PIN vss.gds61
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.982 3.0195 12.042 3.2195 ;
 END
 END vss.gds61
 PIN vss.gds62
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.814 3.0195 11.874 3.2195 ;
 END
 END vss.gds62
 PIN vss.gds63
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 3.0195 13.658 3.2195 ;
 END
 END vss.gds63
 PIN vss.gds64
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 3.0195 11.706 3.2195 ;
 END
 END vss.gds64
 PIN vss.gds65
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.478 3.0195 11.538 3.2195 ;
 END
 END vss.gds65
 PIN vss.gds66
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.31 3.0195 11.37 3.2195 ;
 END
 END vss.gds66
 PIN vss.gds67
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.142 3.0195 11.202 3.2195 ;
 END
 END vss.gds67
 PIN vss.gds68
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.806 3.0195 10.866 3.2195 ;
 END
 END vss.gds68
 PIN vss.gds69
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.638 3.0195 10.698 3.2195 ;
 END
 END vss.gds69
 PIN vss.gds70
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.47 3.0195 10.53 3.2195 ;
 END
 END vss.gds70
 PIN vss.gds71
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 3.0195 11.034 3.2195 ;
 END
 END vss.gds71
 PIN vss.gds72
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 3.06 15.162 3.26 ;
 END
 END vss.gds72
 PIN vss.gds73
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 3.0195 10.362 3.2195 ;
 END
 END vss.gds73
 PIN vss.gds74
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 3.06 14.498 3.26 ;
 END
 END vss.gds74
 PIN vss.gds75
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.262 3.072 13.318 3.272 ;
 END
 END vss.gds75
 PIN vss.gds76
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 2.9235 12.818 3.1235 ;
 END
 END vss.gds76
 PIN vss.gds77
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 2.941 12.378 3.141 ;
 END
 END vss.gds77
 PIN vss.gds78
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 2.803 12.59 3.003 ;
 END
 END vss.gds78
 PIN vss.gds79
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 3.0755 13.058 3.2755 ;
 END
 END vss.gds79
 PIN vss.gds80
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 1.418 13.898 1.618 ;
 END
 END vss.gds80
 PIN vss.gds81
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 14 1.596 14.056 1.769 ;
 RECT 14.168 1.569 14.224 1.769 ;
 RECT 14 2.856 14.056 3.029 ;
 RECT 14.168 2.829 14.224 3.029 ;
 RECT 14 4.116 14.056 4.289 ;
 RECT 14.168 4.089 14.224 4.289 ;
 RECT 14 5.376 14.056 5.549 ;
 RECT 14.168 5.349 14.224 5.549 ;
 RECT 14.336 2.189 14.392 2.389 ;
 RECT 14.168 2.189 14.224 2.389 ;
 RECT 14.336 3.449 14.392 3.649 ;
 RECT 14.168 3.449 14.224 3.649 ;
 RECT 14.336 4.709 14.392 4.909 ;
 RECT 14.168 4.709 14.224 4.909 ;
 RECT 15.008 4.919 15.064 5.119 ;
 RECT 14.84 5.393 14.896 5.558 ;
 RECT 14.672 5.393 14.728 5.558 ;
 RECT 13.664 4.843 13.72 5.043 ;
 RECT 15.008 3.659 15.064 3.859 ;
 RECT 14.84 4.133 14.896 4.298 ;
 RECT 14.672 4.133 14.728 4.298 ;
 RECT 13.664 3.583 13.72 3.783 ;
 RECT 15.008 2.399 15.064 2.599 ;
 RECT 14.84 2.873 14.896 3.038 ;
 RECT 14.672 2.873 14.728 3.038 ;
 RECT 13.664 2.323 13.72 2.523 ;
 RECT 14.336 0.929 14.392 1.129 ;
 RECT 14.168 0.929 14.224 1.129 ;
 RECT 15.008 1.139 15.064 1.339 ;
 RECT 14.84 1.613 14.896 1.778 ;
 RECT 14.672 1.613 14.728 1.778 ;
 RECT 15.176 3.0995 15.232 3.2995 ;
 RECT 13.664 1.063 13.72 1.263 ;
 RECT 12.824 2.884 12.88 3.084 ;
 RECT 13.496 2.895 13.552 3.095 ;
 RECT 13.328 2.833 13.384 3.033 ;
 RECT 13.16 2.884 13.216 3.084 ;
 RECT 12.488 2.914 12.544 3.114 ;
 RECT 12.992 2.884 13.048 3.084 ;
 RECT 12.656 2.914 12.712 3.114 ;
 END
 END vss.gds81
 PIN vss.gds82
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 4.693 16.146 4.893 ;
 END
 END vss.gds82
 PIN vss.gds83
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.986 2.803 18.026 3.003 ;
 END
 END vss.gds83
 PIN vss.gds84
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.206 3.0195 19.266 3.2195 ;
 END
 END vss.gds84
 PIN vss.gds85
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.038 3.0195 19.098 3.2195 ;
 END
 END vss.gds85
 PIN vss.gds86
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.702 3.0195 18.762 3.2195 ;
 END
 END vss.gds86
 PIN vss.gds87
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 3.0195 20.274 3.2195 ;
 END
 END vss.gds87
 PIN vss.gds88
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.374 3.0195 19.434 3.2195 ;
 END
 END vss.gds88
 PIN vss.gds89
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 3.072 16.814 3.272 ;
 END
 END vss.gds89
 PIN vss.gds90
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 2.916 15.418 3.116 ;
 END
 END vss.gds90
 PIN vss.gds91
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 3.0195 19.602 3.2195 ;
 END
 END vss.gds91
 PIN vss.gds92
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 3.0195 18.93 3.2195 ;
 END
 END vss.gds92
 PIN vss.gds93
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 2.9785 16.994 3.1785 ;
 END
 END vss.gds93
 PIN vss.gds94
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 3.06 15.842 3.26 ;
 END
 END vss.gds94
 PIN vss.gds95
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.534 3.0195 18.594 3.2195 ;
 END
 END vss.gds95
 PIN vss.gds96
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.71 3.0195 19.77 3.2195 ;
 END
 END vss.gds96
 PIN vss.gds97
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 3.433 16.146 3.633 ;
 END
 END vss.gds97
 PIN vss.gds98
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.878 3.0195 19.938 3.2195 ;
 END
 END vss.gds98
 PIN vss.gds99
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 2.9235 17.834 3.1235 ;
 END
 END vss.gds99
 PIN vss.gds100
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.438 3.0755 17.494 3.2755 ;
 END
 END vss.gds100
 PIN vss.gds101
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.366 3.0195 18.426 3.2195 ;
 END
 END vss.gds101
 PIN vss.gds102
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.046 3.0195 20.106 3.2195 ;
 END
 END vss.gds102
 PIN vss.gds103
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 2.8265 16.49 3.0265 ;
 END
 END vss.gds103
 PIN vss.gds104
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 2.173 16.146 2.373 ;
 END
 END vss.gds104
 PIN vss.gds105
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 0.913 16.146 1.113 ;
 END
 END vss.gds105
 PIN vss.gds106
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 2.941 18.258 3.141 ;
 END
 END vss.gds106
 PIN vss.gds107
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 2.9235 17.314 3.1235 ;
 END
 END vss.gds107
 PIN vss.gds108
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 15.596 0.58 15.652 0.78 ;
 RECT 15.848 0.583 15.904 0.783 ;
 RECT 16.52 1.616 16.576 1.769 ;
 RECT 15.764 1.613 15.82 1.778 ;
 RECT 15.596 1.613 15.652 1.778 ;
 RECT 15.596 1.84 15.652 2.04 ;
 RECT 15.848 1.843 15.904 2.043 ;
 RECT 16.52 2.876 16.576 3.029 ;
 RECT 15.764 2.873 15.82 3.038 ;
 RECT 15.596 2.873 15.652 3.038 ;
 RECT 15.596 3.1 15.652 3.3 ;
 RECT 15.848 3.103 15.904 3.303 ;
 RECT 16.52 4.136 16.576 4.289 ;
 RECT 15.764 4.133 15.82 4.298 ;
 RECT 15.596 4.133 15.652 4.298 ;
 RECT 15.596 4.36 15.652 4.56 ;
 RECT 15.848 4.363 15.904 4.563 ;
 RECT 16.52 5.396 16.576 5.549 ;
 RECT 15.764 5.393 15.82 5.558 ;
 RECT 15.596 5.393 15.652 5.558 ;
 RECT 15.428 4.919 15.484 5.119 ;
 RECT 16.856 4.7675 16.912 4.9675 ;
 RECT 16.352 5.0195 16.408 5.2195 ;
 RECT 15.428 3.659 15.484 3.859 ;
 RECT 16.352 3.7595 16.408 3.9595 ;
 RECT 16.856 3.5075 16.912 3.7075 ;
 RECT 15.428 2.399 15.484 2.599 ;
 RECT 16.352 2.4995 16.408 2.6995 ;
 RECT 16.856 2.2475 16.912 2.4475 ;
 RECT 15.428 1.139 15.484 1.339 ;
 RECT 16.352 1.2395 16.408 1.4395 ;
 RECT 16.856 0.9875 16.912 1.1875 ;
 RECT 17.864 2.914 17.92 3.114 ;
 RECT 17.696 2.9215 17.752 3.1215 ;
 RECT 17.528 2.914 17.584 3.114 ;
 RECT 17.36 2.914 17.416 3.114 ;
 RECT 17.192 2.914 17.248 3.114 ;
 RECT 17.024 3.029 17.08 3.229 ;
 RECT 18.032 2.914 18.088 3.114 ;
 END
 END vss.gds108
 PIN vss.gds109
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.17 3.0195 25.23 3.2195 ;
 END
 END vss.gds109
 PIN vss.gds110
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.002 3.0195 25.062 3.2195 ;
 END
 END vss.gds110
 PIN vss.gds111
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.834 3.0195 24.894 3.2195 ;
 END
 END vss.gds111
 PIN vss.gds112
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.498 3.0195 24.558 3.2195 ;
 END
 END vss.gds112
 PIN vss.gds113
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.33 3.0195 24.39 3.2195 ;
 END
 END vss.gds113
 PIN vss.gds114
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.162 3.0195 24.222 3.2195 ;
 END
 END vss.gds114
 PIN vss.gds115
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.406 3.0195 23.466 3.2195 ;
 END
 END vss.gds115
 PIN vss.gds116
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.238 3.0195 23.298 3.2195 ;
 END
 END vss.gds116
 PIN vss.gds117
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.07 3.0195 23.13 3.2195 ;
 END
 END vss.gds117
 PIN vss.gds118
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.734 3.0195 22.794 3.2195 ;
 END
 END vss.gds118
 PIN vss.gds119
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.566 3.0195 22.626 3.2195 ;
 END
 END vss.gds119
 PIN vss.gds120
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.398 3.0195 22.458 3.2195 ;
 END
 END vss.gds120
 PIN vss.gds121
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.062 3.0195 22.122 3.2195 ;
 END
 END vss.gds121
 PIN vss.gds122
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.894 3.0195 21.954 3.2195 ;
 END
 END vss.gds122
 PIN vss.gds123
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.726 3.0195 21.786 3.2195 ;
 END
 END vss.gds123
 PIN vss.gds124
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.39 3.0195 21.45 3.2195 ;
 END
 END vss.gds124
 PIN vss.gds125
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.222 3.0195 21.282 3.2195 ;
 END
 END vss.gds125
 PIN vss.gds126
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.054 3.0195 21.114 3.2195 ;
 END
 END vss.gds126
 PIN vss.gds127
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.718 3.0195 20.778 3.2195 ;
 END
 END vss.gds127
 PIN vss.gds128
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.55 3.0195 20.61 3.2195 ;
 END
 END vss.gds128
 PIN vss.gds129
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.382 3.0195 20.442 3.2195 ;
 END
 END vss.gds129
 PIN vss.gds130
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 3.0195 24.726 3.2195 ;
 END
 END vss.gds130
 PIN vss.gds131
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 3.0195 22.962 3.2195 ;
 END
 END vss.gds131
 PIN vss.gds132
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 3.0195 22.29 3.2195 ;
 END
 END vss.gds132
 PIN vss.gds133
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 3.0195 21.618 3.2195 ;
 END
 END vss.gds133
 PIN vss.gds134
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 3.0195 20.946 3.2195 ;
 END
 END vss.gds134
 PIN vss.gds135
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 3.0195 23.634 3.2195 ;
 END
 END vss.gds135
 PIN vss.gds136
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 23.912 4.856 23.968 5.056 ;
 RECT 23.912 3.596 23.968 3.796 ;
 RECT 23.912 2.336 23.968 2.536 ;
 RECT 23.912 1.076 23.968 1.276 ;
 RECT 23.744 2.966 23.8 3.166 ;
 END
 END vss.gds136
 PIN vss.gds137
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.202 3.0195 29.262 3.2195 ;
 END
 END vss.gds137
 PIN vss.gds138
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.034 3.0195 29.094 3.2195 ;
 END
 END vss.gds138
 PIN vss.gds139
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.866 3.0195 28.926 3.2195 ;
 END
 END vss.gds139
 PIN vss.gds140
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.53 3.0195 28.59 3.2195 ;
 END
 END vss.gds140
 PIN vss.gds141
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.362 3.0195 28.422 3.2195 ;
 END
 END vss.gds141
 PIN vss.gds142
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.194 3.0195 28.254 3.2195 ;
 END
 END vss.gds142
 PIN vss.gds143
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.858 3.0195 27.918 3.2195 ;
 END
 END vss.gds143
 PIN vss.gds144
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.69 3.0195 27.75 3.2195 ;
 END
 END vss.gds144
 PIN vss.gds145
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.522 3.0195 27.582 3.2195 ;
 END
 END vss.gds145
 PIN vss.gds146
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.186 3.0195 27.246 3.2195 ;
 END
 END vss.gds146
 PIN vss.gds147
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.018 3.0195 27.078 3.2195 ;
 END
 END vss.gds147
 PIN vss.gds148
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.85 3.0195 26.91 3.2195 ;
 END
 END vss.gds148
 PIN vss.gds149
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.514 3.0195 26.574 3.2195 ;
 END
 END vss.gds149
 PIN vss.gds150
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.346 3.0195 26.406 3.2195 ;
 END
 END vss.gds150
 PIN vss.gds151
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.178 3.0195 26.238 3.2195 ;
 END
 END vss.gds151
 PIN vss.gds152
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.842 3.0195 25.902 3.2195 ;
 END
 END vss.gds152
 PIN vss.gds153
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.674 3.0195 25.734 3.2195 ;
 END
 END vss.gds153
 PIN vss.gds154
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.506 3.0195 25.566 3.2195 ;
 END
 END vss.gds154
 PIN vss.gds155
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 3.0755 30.11 3.2755 ;
 END
 END vss.gds155
 PIN vss.gds156
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 2.941 29.43 3.141 ;
 END
 END vss.gds156
 PIN vss.gds157
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 3.0195 28.758 3.2195 ;
 END
 END vss.gds157
 PIN vss.gds158
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 3.0195 28.086 3.2195 ;
 END
 END vss.gds158
 PIN vss.gds159
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 3.0195 27.414 3.2195 ;
 END
 END vss.gds159
 PIN vss.gds160
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 3.0195 26.742 3.2195 ;
 END
 END vss.gds160
 PIN vss.gds161
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 3.0195 26.07 3.2195 ;
 END
 END vss.gds161
 PIN vss.gds162
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 3.0195 25.398 3.2195 ;
 END
 END vss.gds162
 PIN vss.gds163
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 2.9235 29.87 3.1235 ;
 END
 END vss.gds163
 PIN vss.gds164
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 2.803 29.642 3.003 ;
 END
 END vss.gds164
 PIN vss.gds165
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.876 2.884 29.932 3.084 ;
 RECT 29.54 2.914 29.596 3.114 ;
 RECT 30.212 2.884 30.268 3.084 ;
 RECT 30.044 2.884 30.1 3.084 ;
 RECT 29.708 2.914 29.764 3.114 ;
 END
 END vss.gds165
 PIN vss.gds166
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 1.418 30.95 1.618 ;
 END
 END vss.gds166
 PIN vss.gds167
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 1.458 31.922 1.658 ;
 END
 END vss.gds167
 PIN vss.gds168
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 2.718 31.922 2.918 ;
 END
 END vss.gds168
 PIN vss.gds169
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 3.938 30.95 4.138 ;
 END
 END vss.gds169
 PIN vss.gds170
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 3.978 31.922 4.178 ;
 END
 END vss.gds170
 PIN vss.gds171
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.038 2.803 35.078 3.003 ;
 END
 END vss.gds171
 PIN vss.gds172
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 5.198 30.95 5.398 ;
 END
 END vss.gds172
 PIN vss.gds173
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 5.238 31.922 5.438 ;
 END
 END vss.gds173
 PIN vss.gds174
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.314 3.072 30.37 3.272 ;
 END
 END vss.gds174
 PIN vss.gds175
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 3.06 32.894 3.26 ;
 END
 END vss.gds175
 PIN vss.gds176
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 3.06 32.214 3.26 ;
 END
 END vss.gds176
 PIN vss.gds177
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 2.916 32.47 3.116 ;
 END
 END vss.gds177
 PIN vss.gds178
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 3.0195 30.71 3.2195 ;
 END
 END vss.gds178
 PIN vss.gds179
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 2.8265 33.542 3.0265 ;
 END
 END vss.gds179
 PIN vss.gds180
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 3.06 31.55 3.26 ;
 END
 END vss.gds180
 PIN vss.gds181
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 4.693 33.198 4.893 ;
 END
 END vss.gds181
 PIN vss.gds182
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 2.173 33.198 2.373 ;
 END
 END vss.gds182
 PIN vss.gds183
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 3.072 33.866 3.272 ;
 END
 END vss.gds183
 PIN vss.gds184
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 3.433 33.198 3.633 ;
 END
 END vss.gds184
 PIN vss.gds185
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 2.9235 34.886 3.1235 ;
 END
 END vss.gds185
 PIN vss.gds186
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.49 3.0755 34.546 3.2755 ;
 END
 END vss.gds186
 PIN vss.gds187
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 2.9785 34.046 3.1785 ;
 END
 END vss.gds187
 PIN vss.gds188
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 2.9235 34.366 3.1235 ;
 END
 END vss.gds188
 PIN vss.gds189
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 2.678 30.95 2.878 ;
 END
 END vss.gds189
 PIN vss.gds190
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 0.913 33.198 1.113 ;
 END
 END vss.gds190
 PIN vss.gds191
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 32.648 0.58 32.704 0.78 ;
 RECT 32.9 0.583 32.956 0.783 ;
 RECT 33.572 1.616 33.628 1.769 ;
 RECT 31.052 1.596 31.108 1.769 ;
 RECT 31.22 1.569 31.276 1.769 ;
 RECT 32.816 1.613 32.872 1.778 ;
 RECT 32.648 1.613 32.704 1.778 ;
 RECT 31.892 1.613 31.948 1.778 ;
 RECT 31.724 1.613 31.78 1.778 ;
 RECT 31.388 0.929 31.444 1.129 ;
 RECT 31.22 0.929 31.276 1.129 ;
 RECT 30.716 1.063 30.772 1.263 ;
 RECT 32.648 1.84 32.704 2.04 ;
 RECT 32.9 1.843 32.956 2.043 ;
 RECT 33.572 2.876 33.628 3.029 ;
 RECT 31.052 2.856 31.108 3.029 ;
 RECT 31.22 2.829 31.276 3.029 ;
 RECT 32.816 2.873 32.872 3.038 ;
 RECT 32.648 2.873 32.704 3.038 ;
 RECT 31.892 2.873 31.948 3.038 ;
 RECT 31.724 2.873 31.78 3.038 ;
 RECT 33.572 4.136 33.628 4.289 ;
 RECT 31.052 4.116 31.108 4.289 ;
 RECT 31.22 4.089 31.276 4.289 ;
 RECT 32.816 4.133 32.872 4.298 ;
 RECT 32.648 4.133 32.704 4.298 ;
 RECT 31.892 4.133 31.948 4.298 ;
 RECT 31.724 4.133 31.78 4.298 ;
 RECT 32.648 3.1 32.704 3.3 ;
 RECT 32.9 3.103 32.956 3.303 ;
 RECT 33.572 5.396 33.628 5.549 ;
 RECT 31.052 5.376 31.108 5.549 ;
 RECT 31.22 5.349 31.276 5.549 ;
 RECT 32.816 5.393 32.872 5.558 ;
 RECT 32.648 5.393 32.704 5.558 ;
 RECT 31.892 5.393 31.948 5.558 ;
 RECT 31.724 5.393 31.78 5.558 ;
 RECT 32.648 4.36 32.704 4.56 ;
 RECT 32.9 4.363 32.956 4.563 ;
 RECT 31.388 4.709 31.444 4.909 ;
 RECT 31.22 4.709 31.276 4.909 ;
 RECT 32.06 1.139 32.116 1.339 ;
 RECT 32.48 1.139 32.536 1.339 ;
 RECT 31.388 2.189 31.444 2.389 ;
 RECT 31.22 2.189 31.276 2.389 ;
 RECT 32.06 2.399 32.116 2.599 ;
 RECT 32.48 2.399 32.536 2.599 ;
 RECT 30.716 2.323 30.772 2.523 ;
 RECT 33.404 2.4995 33.46 2.6995 ;
 RECT 33.908 2.2475 33.964 2.4475 ;
 RECT 31.388 3.449 31.444 3.649 ;
 RECT 31.22 3.449 31.276 3.649 ;
 RECT 33.404 3.7595 33.46 3.9595 ;
 RECT 33.908 3.5075 33.964 3.7075 ;
 RECT 30.716 4.843 30.772 5.043 ;
 RECT 32.06 4.919 32.116 5.119 ;
 RECT 32.48 4.919 32.536 5.119 ;
 RECT 30.716 3.583 30.772 3.783 ;
 RECT 32.06 3.659 32.116 3.859 ;
 RECT 32.48 3.659 32.536 3.859 ;
 RECT 30.548 2.895 30.604 3.095 ;
 RECT 33.404 5.0195 33.46 5.2195 ;
 RECT 33.908 4.7675 33.964 4.9675 ;
 RECT 33.404 1.2395 33.46 1.4395 ;
 RECT 33.908 0.9875 33.964 1.1875 ;
 RECT 30.38 2.833 30.436 3.033 ;
 RECT 32.228 3.0995 32.284 3.2995 ;
 RECT 34.916 2.914 34.972 3.114 ;
 RECT 34.748 2.9215 34.804 3.1215 ;
 RECT 34.58 2.914 34.636 3.114 ;
 RECT 34.412 2.914 34.468 3.114 ;
 RECT 34.244 2.914 34.3 3.114 ;
 RECT 35.084 2.914 35.14 3.114 ;
 RECT 34.076 3.029 34.132 3.229 ;
 END
 END vss.gds191
 PIN vss.gds192
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.122 3.0195 40.182 3.2195 ;
 END
 END vss.gds192
 PIN vss.gds193
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.586 3.0195 35.646 3.2195 ;
 END
 END vss.gds193
 PIN vss.gds194
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.754 3.0195 35.814 3.2195 ;
 END
 END vss.gds194
 PIN vss.gds195
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.09 3.0195 36.15 3.2195 ;
 END
 END vss.gds195
 PIN vss.gds196
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.258 3.0195 36.318 3.2195 ;
 END
 END vss.gds196
 PIN vss.gds197
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.426 3.0195 36.486 3.2195 ;
 END
 END vss.gds197
 PIN vss.gds198
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.762 3.0195 36.822 3.2195 ;
 END
 END vss.gds198
 PIN vss.gds199
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.93 3.0195 36.99 3.2195 ;
 END
 END vss.gds199
 PIN vss.gds200
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.098 3.0195 37.158 3.2195 ;
 END
 END vss.gds200
 PIN vss.gds201
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.434 3.0195 37.494 3.2195 ;
 END
 END vss.gds201
 PIN vss.gds202
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.602 3.0195 37.662 3.2195 ;
 END
 END vss.gds202
 PIN vss.gds203
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.77 3.0195 37.83 3.2195 ;
 END
 END vss.gds203
 PIN vss.gds204
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.106 3.0195 38.166 3.2195 ;
 END
 END vss.gds204
 PIN vss.gds205
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.274 3.0195 38.334 3.2195 ;
 END
 END vss.gds205
 PIN vss.gds206
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.442 3.0195 38.502 3.2195 ;
 END
 END vss.gds206
 PIN vss.gds207
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.778 3.0195 38.838 3.2195 ;
 END
 END vss.gds207
 PIN vss.gds208
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.946 3.0195 39.006 3.2195 ;
 END
 END vss.gds208
 PIN vss.gds209
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 3.0195 37.998 3.2195 ;
 END
 END vss.gds209
 PIN vss.gds210
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 3.0195 37.326 3.2195 ;
 END
 END vss.gds210
 PIN vss.gds211
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 3.0195 38.67 3.2195 ;
 END
 END vss.gds211
 PIN vss.gds212
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.45 3.0195 39.51 3.2195 ;
 END
 END vss.gds212
 PIN vss.gds213
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 3.0195 36.654 3.2195 ;
 END
 END vss.gds213
 PIN vss.gds214
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.618 3.0195 39.678 3.2195 ;
 END
 END vss.gds214
 PIN vss.gds215
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.786 3.0195 39.846 3.2195 ;
 END
 END vss.gds215
 PIN vss.gds216
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 3.0195 39.342 3.2195 ;
 END
 END vss.gds216
 PIN vss.gds217
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.114 3.0195 39.174 3.2195 ;
 END
 END vss.gds217
 PIN vss.gds218
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 3.0195 40.014 3.2195 ;
 END
 END vss.gds218
 PIN vss.gds219
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.418 3.0195 35.478 3.2195 ;
 END
 END vss.gds219
 PIN vss.gds220
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 2.941 35.31 3.141 ;
 END
 END vss.gds220
 PIN vss.gds221
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 3.0195 35.982 3.2195 ;
 END
 END vss.gds221
 PIN vss.gds222
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.91 3.0195 44.97 3.2195 ;
 END
 END vss.gds222
 PIN vss.gds223
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.742 3.0195 44.802 3.2195 ;
 END
 END vss.gds223
 PIN vss.gds224
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.574 3.0195 44.634 3.2195 ;
 END
 END vss.gds224
 PIN vss.gds225
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.238 3.0195 44.298 3.2195 ;
 END
 END vss.gds225
 PIN vss.gds226
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.07 3.0195 44.13 3.2195 ;
 END
 END vss.gds226
 PIN vss.gds227
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.902 3.0195 43.962 3.2195 ;
 END
 END vss.gds227
 PIN vss.gds228
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.566 3.0195 43.626 3.2195 ;
 END
 END vss.gds228
 PIN vss.gds229
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.398 3.0195 43.458 3.2195 ;
 END
 END vss.gds229
 PIN vss.gds230
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.23 3.0195 43.29 3.2195 ;
 END
 END vss.gds230
 PIN vss.gds231
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.894 3.0195 42.954 3.2195 ;
 END
 END vss.gds231
 PIN vss.gds232
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.726 3.0195 42.786 3.2195 ;
 END
 END vss.gds232
 PIN vss.gds233
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.558 3.0195 42.618 3.2195 ;
 END
 END vss.gds233
 PIN vss.gds234
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.222 3.0195 42.282 3.2195 ;
 END
 END vss.gds234
 PIN vss.gds235
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.054 3.0195 42.114 3.2195 ;
 END
 END vss.gds235
 PIN vss.gds236
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.886 3.0195 41.946 3.2195 ;
 END
 END vss.gds236
 PIN vss.gds237
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.55 3.0195 41.61 3.2195 ;
 END
 END vss.gds237
 PIN vss.gds238
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.382 3.0195 41.442 3.2195 ;
 END
 END vss.gds238
 PIN vss.gds239
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.214 3.0195 41.274 3.2195 ;
 END
 END vss.gds239
 PIN vss.gds240
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.29 3.0195 40.35 3.2195 ;
 END
 END vss.gds240
 PIN vss.gds241
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.458 3.0195 40.518 3.2195 ;
 END
 END vss.gds241
 PIN vss.gds242
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 3.0195 45.138 3.2195 ;
 END
 END vss.gds242
 PIN vss.gds243
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 3.0195 44.466 3.2195 ;
 END
 END vss.gds243
 PIN vss.gds244
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 3.0195 43.794 3.2195 ;
 END
 END vss.gds244
 PIN vss.gds245
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 3.0195 43.122 3.2195 ;
 END
 END vss.gds245
 PIN vss.gds246
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 3.0195 42.45 3.2195 ;
 END
 END vss.gds246
 PIN vss.gds247
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 3.0195 41.778 3.2195 ;
 END
 END vss.gds247
 PIN vss.gds248
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 3.0195 40.686 3.2195 ;
 END
 END vss.gds248
 PIN vss.gds249
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 40.964 4.856 41.02 5.056 ;
 RECT 40.964 3.596 41.02 3.796 ;
 RECT 40.964 2.336 41.02 2.536 ;
 RECT 40.964 1.076 41.02 1.276 ;
 RECT 40.796 2.966 40.852 3.166 ;
 END
 END vss.gds249
 PIN vss.gds250
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 2.173 50.25 2.373 ;
 END
 END vss.gds250
 PIN vss.gds251
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 1.418 48.002 1.618 ;
 END
 END vss.gds251
 PIN vss.gds252
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 1.458 48.974 1.658 ;
 END
 END vss.gds252
 PIN vss.gds253
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 2.718 48.974 2.918 ;
 END
 END vss.gds253
 PIN vss.gds254
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 3.978 48.974 4.178 ;
 END
 END vss.gds254
 PIN vss.gds255
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 2.678 48.002 2.878 ;
 END
 END vss.gds255
 PIN vss.gds256
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 5.198 48.002 5.398 ;
 END
 END vss.gds256
 PIN vss.gds257
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 5.238 48.974 5.438 ;
 END
 END vss.gds257
 PIN vss.gds258
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.366 3.072 47.422 3.272 ;
 END
 END vss.gds258
 PIN vss.gds259
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.254 3.0195 46.314 3.2195 ;
 END
 END vss.gds259
 PIN vss.gds260
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.086 3.0195 46.146 3.2195 ;
 END
 END vss.gds260
 PIN vss.gds261
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.918 3.0195 45.978 3.2195 ;
 END
 END vss.gds261
 PIN vss.gds262
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.582 3.0195 45.642 3.2195 ;
 END
 END vss.gds262
 PIN vss.gds263
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.414 3.0195 45.474 3.2195 ;
 END
 END vss.gds263
 PIN vss.gds264
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.246 3.0195 45.306 3.2195 ;
 END
 END vss.gds264
 PIN vss.gds265
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 3.0195 45.81 3.2195 ;
 END
 END vss.gds265
 PIN vss.gds266
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 2.941 46.482 3.141 ;
 END
 END vss.gds266
 PIN vss.gds267
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 3.0755 47.162 3.2755 ;
 END
 END vss.gds267
 PIN vss.gds268
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 2.9235 46.922 3.1235 ;
 END
 END vss.gds268
 PIN vss.gds269
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 2.803 46.694 3.003 ;
 END
 END vss.gds269
 PIN vss.gds270
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 3.0195 47.762 3.2195 ;
 END
 END vss.gds270
 PIN vss.gds271
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 3.06 49.266 3.26 ;
 END
 END vss.gds271
 PIN vss.gds272
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 4.693 50.25 4.893 ;
 END
 END vss.gds272
 PIN vss.gds273
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 3.433 50.25 3.633 ;
 END
 END vss.gds273
 PIN vss.gds274
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 3.06 48.602 3.26 ;
 END
 END vss.gds274
 PIN vss.gds275
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 3.06 49.946 3.26 ;
 END
 END vss.gds275
 PIN vss.gds276
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 2.916 49.522 3.116 ;
 END
 END vss.gds276
 PIN vss.gds277
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 3.938 48.002 4.138 ;
 END
 END vss.gds277
 PIN vss.gds278
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 0.913 50.25 1.113 ;
 END
 END vss.gds278
 PIN vss.gds279
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 49.7 0.58 49.756 0.78 ;
 RECT 49.952 0.583 50.008 0.783 ;
 RECT 48.104 1.596 48.16 1.769 ;
 RECT 48.272 1.569 48.328 1.769 ;
 RECT 49.868 1.613 49.924 1.778 ;
 RECT 49.7 1.613 49.756 1.778 ;
 RECT 48.944 1.613 49 1.778 ;
 RECT 48.776 1.613 48.832 1.778 ;
 RECT 48.44 0.929 48.496 1.129 ;
 RECT 48.272 0.929 48.328 1.129 ;
 RECT 47.768 1.063 47.824 1.263 ;
 RECT 49.7 4.36 49.756 4.56 ;
 RECT 49.952 4.363 50.008 4.563 ;
 RECT 48.104 2.856 48.16 3.029 ;
 RECT 48.272 2.829 48.328 3.029 ;
 RECT 49.868 2.873 49.924 3.038 ;
 RECT 49.7 2.873 49.756 3.038 ;
 RECT 48.944 2.873 49 3.038 ;
 RECT 48.776 2.873 48.832 3.038 ;
 RECT 48.104 4.116 48.16 4.289 ;
 RECT 48.272 4.089 48.328 4.289 ;
 RECT 49.868 4.133 49.924 4.298 ;
 RECT 49.7 4.133 49.756 4.298 ;
 RECT 48.944 4.133 49 4.298 ;
 RECT 48.776 4.133 48.832 4.298 ;
 RECT 48.104 5.376 48.16 5.549 ;
 RECT 48.272 5.349 48.328 5.549 ;
 RECT 49.868 5.393 49.924 5.558 ;
 RECT 49.7 5.393 49.756 5.558 ;
 RECT 48.944 5.393 49 5.558 ;
 RECT 48.776 5.393 48.832 5.558 ;
 RECT 49.7 3.1 49.756 3.3 ;
 RECT 49.952 3.103 50.008 3.303 ;
 RECT 49.7 1.84 49.756 2.04 ;
 RECT 49.952 1.843 50.008 2.043 ;
 RECT 49.112 1.139 49.168 1.339 ;
 RECT 49.532 1.139 49.588 1.339 ;
 RECT 48.44 4.709 48.496 4.909 ;
 RECT 48.272 4.709 48.328 4.909 ;
 RECT 47.768 4.843 47.824 5.043 ;
 RECT 49.112 4.919 49.168 5.119 ;
 RECT 49.532 4.919 49.588 5.119 ;
 RECT 48.44 3.449 48.496 3.649 ;
 RECT 48.272 3.449 48.328 3.649 ;
 RECT 49.112 3.659 49.168 3.859 ;
 RECT 49.532 3.659 49.588 3.859 ;
 RECT 49.112 2.399 49.168 2.599 ;
 RECT 49.532 2.399 49.588 2.599 ;
 RECT 48.44 2.189 48.496 2.389 ;
 RECT 48.272 2.189 48.328 2.389 ;
 RECT 47.768 2.323 47.824 2.523 ;
 RECT 47.768 3.583 47.824 3.783 ;
 RECT 47.6 2.895 47.656 3.095 ;
 RECT 47.432 2.833 47.488 3.033 ;
 RECT 47.264 2.884 47.32 3.084 ;
 RECT 46.928 2.884 46.984 3.084 ;
 RECT 46.592 2.914 46.648 3.114 ;
 RECT 47.096 2.884 47.152 3.084 ;
 RECT 49.28 3.0995 49.336 3.2995 ;
 RECT 46.76 2.914 46.816 3.114 ;
 END
 END vss.gds279
 PIN vss.gds280
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.09 2.803 52.13 3.003 ;
 END
 END vss.gds280
 PIN vss.gds281
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.638 3.0195 52.698 3.2195 ;
 END
 END vss.gds281
 PIN vss.gds282
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.806 3.0195 52.866 3.2195 ;
 END
 END vss.gds282
 PIN vss.gds283
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.142 3.0195 53.202 3.2195 ;
 END
 END vss.gds283
 PIN vss.gds284
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.31 3.0195 53.37 3.2195 ;
 END
 END vss.gds284
 PIN vss.gds285
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.478 3.0195 53.538 3.2195 ;
 END
 END vss.gds285
 PIN vss.gds286
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.814 3.0195 53.874 3.2195 ;
 END
 END vss.gds286
 PIN vss.gds287
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.982 3.0195 54.042 3.2195 ;
 END
 END vss.gds287
 PIN vss.gds288
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.15 3.0195 54.21 3.2195 ;
 END
 END vss.gds288
 PIN vss.gds289
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.486 3.0195 54.546 3.2195 ;
 END
 END vss.gds289
 PIN vss.gds290
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.654 3.0195 54.714 3.2195 ;
 END
 END vss.gds290
 PIN vss.gds291
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.822 3.0195 54.882 3.2195 ;
 END
 END vss.gds291
 PIN vss.gds292
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.158 3.0195 55.218 3.2195 ;
 END
 END vss.gds292
 PIN vss.gds293
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 3.0195 54.378 3.2195 ;
 END
 END vss.gds293
 PIN vss.gds294
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 3.0195 55.05 3.2195 ;
 END
 END vss.gds294
 PIN vss.gds295
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 3.0195 53.706 3.2195 ;
 END
 END vss.gds295
 PIN vss.gds296
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 2.9235 51.418 3.1235 ;
 END
 END vss.gds296
 PIN vss.gds297
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 3.072 50.918 3.272 ;
 END
 END vss.gds297
 PIN vss.gds298
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 3.0195 53.034 3.2195 ;
 END
 END vss.gds298
 PIN vss.gds299
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 2.9235 51.938 3.1235 ;
 END
 END vss.gds299
 PIN vss.gds300
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 2.8265 50.594 3.0265 ;
 END
 END vss.gds300
 PIN vss.gds301
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.47 3.0195 52.53 3.2195 ;
 END
 END vss.gds301
 PIN vss.gds302
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.542 3.0755 51.598 3.2755 ;
 END
 END vss.gds302
 PIN vss.gds303
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 2.941 52.362 3.141 ;
 END
 END vss.gds303
 PIN vss.gds304
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 2.9785 51.098 3.1785 ;
 END
 END vss.gds304
 PIN vss.gds305
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 50.624 1.616 50.68 1.769 ;
 RECT 50.624 2.876 50.68 3.029 ;
 RECT 50.624 4.136 50.68 4.289 ;
 RECT 50.624 5.396 50.68 5.549 ;
 RECT 50.96 4.7675 51.016 4.9675 ;
 RECT 50.456 5.0195 50.512 5.2195 ;
 RECT 50.456 3.7595 50.512 3.9595 ;
 RECT 50.96 3.5075 51.016 3.7075 ;
 RECT 50.96 2.2475 51.016 2.4475 ;
 RECT 50.456 2.4995 50.512 2.6995 ;
 RECT 50.456 1.2395 50.512 1.4395 ;
 RECT 50.96 0.9875 51.016 1.1875 ;
 RECT 51.968 2.914 52.024 3.114 ;
 RECT 51.8 2.9215 51.856 3.1215 ;
 RECT 51.632 2.914 51.688 3.114 ;
 RECT 51.464 2.914 51.52 3.114 ;
 RECT 51.296 2.914 51.352 3.114 ;
 RECT 52.136 2.914 52.192 3.114 ;
 RECT 51.128 3.029 51.184 3.229 ;
 END
 END vss.gds305
 PIN vss.gds306
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.946 3.0195 60.006 3.2195 ;
 END
 END vss.gds306
 PIN vss.gds307
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.778 3.0195 59.838 3.2195 ;
 END
 END vss.gds307
 PIN vss.gds308
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.61 3.0195 59.67 3.2195 ;
 END
 END vss.gds308
 PIN vss.gds309
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.274 3.0195 59.334 3.2195 ;
 END
 END vss.gds309
 PIN vss.gds310
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.106 3.0195 59.166 3.2195 ;
 END
 END vss.gds310
 PIN vss.gds311
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.938 3.0195 58.998 3.2195 ;
 END
 END vss.gds311
 PIN vss.gds312
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.602 3.0195 58.662 3.2195 ;
 END
 END vss.gds312
 PIN vss.gds313
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.434 3.0195 58.494 3.2195 ;
 END
 END vss.gds313
 PIN vss.gds314
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.266 3.0195 58.326 3.2195 ;
 END
 END vss.gds314
 PIN vss.gds315
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.326 3.0195 55.386 3.2195 ;
 END
 END vss.gds315
 PIN vss.gds316
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.494 3.0195 55.554 3.2195 ;
 END
 END vss.gds316
 PIN vss.gds317
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.83 3.0195 55.89 3.2195 ;
 END
 END vss.gds317
 PIN vss.gds318
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.998 3.0195 56.058 3.2195 ;
 END
 END vss.gds318
 PIN vss.gds319
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.166 3.0195 56.226 3.2195 ;
 END
 END vss.gds319
 PIN vss.gds320
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 3.0195 60.174 3.2195 ;
 END
 END vss.gds320
 PIN vss.gds321
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 3.0195 59.502 3.2195 ;
 END
 END vss.gds321
 PIN vss.gds322
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 3.0195 58.83 3.2195 ;
 END
 END vss.gds322
 PIN vss.gds323
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 3.0195 55.722 3.2195 ;
 END
 END vss.gds323
 PIN vss.gds324
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 3.0195 56.394 3.2195 ;
 END
 END vss.gds324
 PIN vss.gds325
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.502 3.0195 56.562 3.2195 ;
 END
 END vss.gds325
 PIN vss.gds326
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.67 3.0195 56.73 3.2195 ;
 END
 END vss.gds326
 PIN vss.gds327
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.838 3.0195 56.898 3.2195 ;
 END
 END vss.gds327
 PIN vss.gds328
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.342 3.0195 57.402 3.2195 ;
 END
 END vss.gds328
 PIN vss.gds329
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.51 3.0195 57.57 3.2195 ;
 END
 END vss.gds329
 PIN vss.gds330
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 3.0195 57.738 3.2195 ;
 END
 END vss.gds330
 PIN vss.gds331
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 3.0195 57.066 3.2195 ;
 END
 END vss.gds331
 PIN vss.gds332
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.174 3.0195 57.234 3.2195 ;
 END
 END vss.gds332
 PIN vss.gds333
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 58.016 4.856 58.072 5.056 ;
 RECT 58.016 3.596 58.072 3.796 ;
 RECT 58.016 2.336 58.072 2.536 ;
 RECT 58.016 1.076 58.072 1.276 ;
 RECT 57.848 2.966 57.904 3.166 ;
 END
 END vss.gds333
 PIN vss.gds334
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 1.418 65.054 1.618 ;
 END
 END vss.gds334
 PIN vss.gds335
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 3.938 65.054 4.138 ;
 END
 END vss.gds335
 PIN vss.gds336
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 2.678 65.054 2.878 ;
 END
 END vss.gds336
 PIN vss.gds337
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 5.198 65.054 5.398 ;
 END
 END vss.gds337
 PIN vss.gds338
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.418 3.072 64.474 3.272 ;
 END
 END vss.gds338
 PIN vss.gds339
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.306 3.0195 63.366 3.2195 ;
 END
 END vss.gds339
 PIN vss.gds340
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.138 3.0195 63.198 3.2195 ;
 END
 END vss.gds340
 PIN vss.gds341
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.97 3.0195 63.03 3.2195 ;
 END
 END vss.gds341
 PIN vss.gds342
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.634 3.0195 62.694 3.2195 ;
 END
 END vss.gds342
 PIN vss.gds343
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.466 3.0195 62.526 3.2195 ;
 END
 END vss.gds343
 PIN vss.gds344
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.298 3.0195 62.358 3.2195 ;
 END
 END vss.gds344
 PIN vss.gds345
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.962 3.0195 62.022 3.2195 ;
 END
 END vss.gds345
 PIN vss.gds346
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.794 3.0195 61.854 3.2195 ;
 END
 END vss.gds346
 PIN vss.gds347
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.626 3.0195 61.686 3.2195 ;
 END
 END vss.gds347
 PIN vss.gds348
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.29 3.0195 61.35 3.2195 ;
 END
 END vss.gds348
 PIN vss.gds349
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.122 3.0195 61.182 3.2195 ;
 END
 END vss.gds349
 PIN vss.gds350
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.954 3.0195 61.014 3.2195 ;
 END
 END vss.gds350
 PIN vss.gds351
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.618 3.0195 60.678 3.2195 ;
 END
 END vss.gds351
 PIN vss.gds352
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.45 3.0195 60.51 3.2195 ;
 END
 END vss.gds352
 PIN vss.gds353
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.282 3.0195 60.342 3.2195 ;
 END
 END vss.gds353
 PIN vss.gds354
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 3.0755 64.214 3.2755 ;
 END
 END vss.gds354
 PIN vss.gds355
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 2.941 63.534 3.141 ;
 END
 END vss.gds355
 PIN vss.gds356
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 3.0195 62.862 3.2195 ;
 END
 END vss.gds356
 PIN vss.gds357
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 3.0195 62.19 3.2195 ;
 END
 END vss.gds357
 PIN vss.gds358
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 3.0195 61.518 3.2195 ;
 END
 END vss.gds358
 PIN vss.gds359
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 3.0195 60.846 3.2195 ;
 END
 END vss.gds359
 PIN vss.gds360
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 2.9235 63.974 3.1235 ;
 END
 END vss.gds360
 PIN vss.gds361
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 2.803 63.746 3.003 ;
 END
 END vss.gds361
 PIN vss.gds362
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 3.0195 64.814 3.2195 ;
 END
 END vss.gds362
 PIN vss.gds363
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 65.156 1.596 65.212 1.769 ;
 RECT 65.156 2.856 65.212 3.029 ;
 RECT 65.156 4.116 65.212 4.289 ;
 RECT 65.156 5.376 65.212 5.549 ;
 RECT 64.82 1.063 64.876 1.263 ;
 RECT 64.82 4.843 64.876 5.043 ;
 RECT 64.82 2.323 64.876 2.523 ;
 RECT 64.82 3.583 64.876 3.783 ;
 RECT 64.652 2.895 64.708 3.095 ;
 RECT 64.484 2.833 64.54 3.033 ;
 RECT 63.98 2.884 64.036 3.084 ;
 RECT 64.316 2.884 64.372 3.084 ;
 RECT 64.148 2.884 64.204 3.084 ;
 RECT 63.644 2.914 63.7 3.114 ;
 RECT 63.812 2.914 63.868 3.114 ;
 END
 END vss.gds363
 PIN vss.gds364
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 1.458 66.026 1.658 ;
 END
 END vss.gds364
 PIN vss.gds365
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 2.718 66.026 2.918 ;
 END
 END vss.gds365
 PIN vss.gds366
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 3.978 66.026 4.178 ;
 END
 END vss.gds366
 PIN vss.gds367
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 5.238 66.026 5.438 ;
 END
 END vss.gds367
 PIN vss.gds368
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.142 2.803 69.182 3.003 ;
 END
 END vss.gds368
 PIN vss.gds369
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.69 3.0195 69.75 3.2195 ;
 END
 END vss.gds369
 PIN vss.gds370
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.858 3.0195 69.918 3.2195 ;
 END
 END vss.gds370
 PIN vss.gds371
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.194 3.0195 70.254 3.2195 ;
 END
 END vss.gds371
 PIN vss.gds372
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 2.916 66.574 3.116 ;
 END
 END vss.gds372
 PIN vss.gds373
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 3.06 66.318 3.26 ;
 END
 END vss.gds373
 PIN vss.gds374
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 3.0195 70.086 3.2195 ;
 END
 END vss.gds374
 PIN vss.gds375
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 2.9785 68.15 3.1785 ;
 END
 END vss.gds375
 PIN vss.gds376
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 2.8265 67.646 3.0265 ;
 END
 END vss.gds376
 PIN vss.gds377
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 3.072 67.97 3.272 ;
 END
 END vss.gds377
 PIN vss.gds378
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 3.06 65.654 3.26 ;
 END
 END vss.gds378
 PIN vss.gds379
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 3.06 66.998 3.26 ;
 END
 END vss.gds379
 PIN vss.gds380
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 2.9235 68.99 3.1235 ;
 END
 END vss.gds380
 PIN vss.gds381
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 4.693 67.302 4.893 ;
 END
 END vss.gds381
 PIN vss.gds382
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 3.433 67.302 3.633 ;
 END
 END vss.gds382
 PIN vss.gds383
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.594 3.0755 68.65 3.2755 ;
 END
 END vss.gds383
 PIN vss.gds384
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 2.9235 68.47 3.1235 ;
 END
 END vss.gds384
 PIN vss.gds385
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 2.173 67.302 2.373 ;
 END
 END vss.gds385
 PIN vss.gds386
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 0.913 67.302 1.113 ;
 END
 END vss.gds386
 PIN vss.gds387
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.522 3.0195 69.582 3.2195 ;
 END
 END vss.gds387
 PIN vss.gds388
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 2.941 69.414 3.141 ;
 END
 END vss.gds388
 PIN vss.gds389
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 67.676 1.616 67.732 1.769 ;
 RECT 65.324 1.569 65.38 1.769 ;
 RECT 66.92 1.613 66.976 1.778 ;
 RECT 66.752 1.613 66.808 1.778 ;
 RECT 65.996 1.613 66.052 1.778 ;
 RECT 65.828 1.613 65.884 1.778 ;
 RECT 66.752 0.58 66.808 0.78 ;
 RECT 67.004 0.583 67.06 0.783 ;
 RECT 67.676 2.876 67.732 3.029 ;
 RECT 65.324 2.829 65.38 3.029 ;
 RECT 66.92 2.873 66.976 3.038 ;
 RECT 66.752 2.873 66.808 3.038 ;
 RECT 65.996 2.873 66.052 3.038 ;
 RECT 65.828 2.873 65.884 3.038 ;
 RECT 67.676 4.136 67.732 4.289 ;
 RECT 65.324 4.089 65.38 4.289 ;
 RECT 66.92 4.133 66.976 4.298 ;
 RECT 66.752 4.133 66.808 4.298 ;
 RECT 65.996 4.133 66.052 4.298 ;
 RECT 65.828 4.133 65.884 4.298 ;
 RECT 67.676 5.396 67.732 5.549 ;
 RECT 65.324 5.349 65.38 5.549 ;
 RECT 66.92 5.393 66.976 5.558 ;
 RECT 66.752 5.393 66.808 5.558 ;
 RECT 65.996 5.393 66.052 5.558 ;
 RECT 65.828 5.393 65.884 5.558 ;
 RECT 65.492 0.929 65.548 1.129 ;
 RECT 65.324 0.929 65.38 1.129 ;
 RECT 66.752 3.1 66.808 3.3 ;
 RECT 67.004 3.103 67.06 3.303 ;
 RECT 66.752 1.84 66.808 2.04 ;
 RECT 67.004 1.843 67.06 2.043 ;
 RECT 65.492 2.189 65.548 2.389 ;
 RECT 65.324 2.189 65.38 2.389 ;
 RECT 66.752 4.36 66.808 4.56 ;
 RECT 67.004 4.363 67.06 4.563 ;
 RECT 66.164 1.139 66.22 1.339 ;
 RECT 66.584 1.139 66.64 1.339 ;
 RECT 67.508 5.0195 67.564 5.2195 ;
 RECT 68.012 4.7675 68.068 4.9675 ;
 RECT 65.492 4.709 65.548 4.909 ;
 RECT 65.324 4.709 65.38 4.909 ;
 RECT 66.164 4.919 66.22 5.119 ;
 RECT 66.584 4.919 66.64 5.119 ;
 RECT 66.164 2.399 66.22 2.599 ;
 RECT 66.584 2.399 66.64 2.599 ;
 RECT 68.012 3.5075 68.068 3.7075 ;
 RECT 67.508 3.7595 67.564 3.9595 ;
 RECT 66.164 3.659 66.22 3.859 ;
 RECT 66.584 3.659 66.64 3.859 ;
 RECT 65.492 3.449 65.548 3.649 ;
 RECT 65.324 3.449 65.38 3.649 ;
 RECT 67.508 2.4995 67.564 2.6995 ;
 RECT 68.012 2.2475 68.068 2.4475 ;
 RECT 66.332 3.0995 66.388 3.2995 ;
 RECT 67.508 1.2395 67.564 1.4395 ;
 RECT 68.012 0.9875 68.068 1.1875 ;
 RECT 69.02 2.914 69.076 3.114 ;
 RECT 68.852 2.9215 68.908 3.1215 ;
 RECT 68.684 2.914 68.74 3.114 ;
 RECT 68.516 2.914 68.572 3.114 ;
 RECT 68.348 2.914 68.404 3.114 ;
 RECT 69.188 2.914 69.244 3.114 ;
 RECT 68.18 3.029 68.236 3.229 ;
 END
 END vss.gds389
 PIN vss.gds390
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.362 3.0195 70.422 3.2195 ;
 END
 END vss.gds390
 PIN vss.gds391
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.53 3.0195 70.59 3.2195 ;
 END
 END vss.gds391
 PIN vss.gds392
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.866 3.0195 70.926 3.2195 ;
 END
 END vss.gds392
 PIN vss.gds393
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.034 3.0195 71.094 3.2195 ;
 END
 END vss.gds393
 PIN vss.gds394
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.202 3.0195 71.262 3.2195 ;
 END
 END vss.gds394
 PIN vss.gds395
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.538 3.0195 71.598 3.2195 ;
 END
 END vss.gds395
 PIN vss.gds396
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.706 3.0195 71.766 3.2195 ;
 END
 END vss.gds396
 PIN vss.gds397
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.874 3.0195 71.934 3.2195 ;
 END
 END vss.gds397
 PIN vss.gds398
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.21 3.0195 72.27 3.2195 ;
 END
 END vss.gds398
 PIN vss.gds399
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.378 3.0195 72.438 3.2195 ;
 END
 END vss.gds399
 PIN vss.gds400
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.546 3.0195 72.606 3.2195 ;
 END
 END vss.gds400
 PIN vss.gds401
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.882 3.0195 72.942 3.2195 ;
 END
 END vss.gds401
 PIN vss.gds402
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.05 3.0195 73.11 3.2195 ;
 END
 END vss.gds402
 PIN vss.gds403
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 3.0195 71.43 3.2195 ;
 END
 END vss.gds403
 PIN vss.gds404
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 3.0195 72.102 3.2195 ;
 END
 END vss.gds404
 PIN vss.gds405
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 3.0195 72.774 3.2195 ;
 END
 END vss.gds405
 PIN vss.gds406
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 3.0195 70.758 3.2195 ;
 END
 END vss.gds406
 PIN vss.gds407
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.554 3.0195 73.614 3.2195 ;
 END
 END vss.gds407
 PIN vss.gds408
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.722 3.0195 73.782 3.2195 ;
 END
 END vss.gds408
 PIN vss.gds409
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.89 3.0195 73.95 3.2195 ;
 END
 END vss.gds409
 PIN vss.gds410
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 3.0195 74.118 3.2195 ;
 END
 END vss.gds410
 PIN vss.gds411
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.394 3.0195 74.454 3.2195 ;
 END
 END vss.gds411
 PIN vss.gds412
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.562 3.0195 74.622 3.2195 ;
 END
 END vss.gds412
 PIN vss.gds413
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 3.0195 74.79 3.2195 ;
 END
 END vss.gds413
 PIN vss.gds414
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.218 3.0195 73.278 3.2195 ;
 END
 END vss.gds414
 PIN vss.gds415
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 3.0195 73.446 3.2195 ;
 END
 END vss.gds415
 PIN vss.gds416
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.226 3.0195 74.286 3.2195 ;
 END
 END vss.gds416
 PIN vss.gds417
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 7.6805 0.29 7.8805 ;
 END
 END vss.gds417
 PIN vss.gds418
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 5.953 2.962 6.153 ;
 END
 END vss.gds418
 PIN vss.gds419
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 9.733 2.962 9.933 ;
 END
 END vss.gds419
 PIN vss.gds420
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 6.812 3.142 7.012 ;
 END
 END vss.gds420
 PIN vss.gds421
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 5.552 3.142 5.752 ;
 END
 END vss.gds421
 PIN vss.gds422
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 8.473 2.962 8.673 ;
 END
 END vss.gds422
 PIN vss.gds423
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 8.072 3.142 8.272 ;
 END
 END vss.gds423
 PIN vss.gds424
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 7.213 2.962 7.413 ;
 END
 END vss.gds424
 PIN vss.gds425
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.286 7.843 3.326 8.043 ;
 END
 END vss.gds425
 PIN vss.gds426
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.754 7.843 3.794 8.043 ;
 END
 END vss.gds426
 PIN vss.gds427
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.442 7.437 4.482 7.637 ;
 END
 END vss.gds427
 PIN vss.gds428
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 9.332 3.142 9.532 ;
 END
 END vss.gds428
 PIN vss.gds429
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 7.638 0.602 7.838 ;
 END
 END vss.gds429
 PIN vss.gds430
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.414 8.119 3.454 8.319 ;
 END
 END vss.gds430
 PIN vss.gds431
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 7.437 0.942 7.637 ;
 END
 END vss.gds431
 PIN vss.gds432
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 7.981 1.282 8.181 ;
 END
 END vss.gds432
 PIN vss.gds433
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 7.8665 2.122 8.0665 ;
 END
 END vss.gds433
 PIN vss.gds434
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 7.437 4.882 7.637 ;
 END
 END vss.gds434
 PIN vss.gds435
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.57 7.64 4.61 7.84 ;
 END
 END vss.gds435
 PIN vss.gds436
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 8.831 4.194 9.031 ;
 END
 END vss.gds436
 PIN vss.gds437
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 7.843 5.074 8.043 ;
 END
 END vss.gds437
 PIN vss.gds438
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.562 8.119 3.602 8.319 ;
 END
 END vss.gds438
 PIN vss.gds439
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 7.7395 4.002 7.9395 ;
 END
 END vss.gds439
 PIN vss.gds440
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 7.7395 5.282 7.9395 ;
 END
 END vss.gds440
 PIN vss.gds441
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 7.778 2.302 7.978 ;
 END
 END vss.gds441
 PIN vss.gds442
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 8.2155 1.462 8.4155 ;
 END
 END vss.gds442
 PIN vss.gds443
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 7.5375 0.718 7.7375 ;
 END
 END vss.gds443
 PIN vss.gds444
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 2.576 5.9535 2.632 6.1535 ;
 RECT 2.408 5.9535 2.464 6.1535 ;
 RECT 2.996 5.9535 3.052 6.1535 ;
 RECT 3.332 6.045 3.388 6.245 ;
 RECT 3.5 6.0015 3.556 6.2015 ;
 RECT 0.98 5.8685 1.036 6.0685 ;
 RECT 2.072 5.869 2.128 6.069 ;
 RECT 2.576 7.2135 2.632 7.4135 ;
 RECT 2.408 7.2135 2.464 7.4135 ;
 RECT 2.996 7.2135 3.052 7.4135 ;
 RECT 3.332 7.305 3.388 7.505 ;
 RECT 3.5 7.2615 3.556 7.4615 ;
 RECT 0.98 7.1285 1.036 7.3285 ;
 RECT 2.072 7.129 2.128 7.329 ;
 RECT 2.576 8.4735 2.632 8.6735 ;
 RECT 2.408 8.4735 2.464 8.6735 ;
 RECT 2.996 8.4735 3.052 8.6735 ;
 RECT 3.332 8.565 3.388 8.765 ;
 RECT 3.5 8.5215 3.556 8.7215 ;
 RECT 0.98 8.3885 1.036 8.5885 ;
 RECT 2.072 8.389 2.128 8.589 ;
 RECT 2.576 9.7335 2.632 9.9335 ;
 RECT 2.408 9.7335 2.464 9.9335 ;
 RECT 2.996 9.7335 3.052 9.9335 ;
 RECT 3.332 9.825 3.388 10.025 ;
 RECT 3.5 9.7815 3.556 9.9815 ;
 RECT 0.98 9.6485 1.036 9.8485 ;
 RECT 2.072 9.649 2.128 9.849 ;
 RECT 0.392 9.739 0.448 9.939 ;
 RECT 0.812 9.825 0.868 10.025 ;
 RECT 0.644 9.739 0.7 9.939 ;
 RECT 1.232 9.739 1.288 9.939 ;
 RECT 1.4 9.739 1.456 9.939 ;
 RECT 1.568 9.739 1.624 9.939 ;
 RECT 1.82 9.739 1.876 9.939 ;
 RECT 2.24 9.739 2.296 9.939 ;
 RECT 2.744 9.649 2.8 9.849 ;
 RECT 3.164 9.739 3.22 9.939 ;
 RECT 3.92 9.739 3.976 9.939 ;
 RECT 3.752 10.009 3.808 10.209 ;
 RECT 4.508 9.9385 4.564 10.1385 ;
 RECT 0.392 8.479 0.448 8.679 ;
 RECT 0.812 8.565 0.868 8.765 ;
 RECT 0.644 8.479 0.7 8.679 ;
 RECT 1.232 8.479 1.288 8.679 ;
 RECT 1.4 8.479 1.456 8.679 ;
 RECT 1.568 8.479 1.624 8.679 ;
 RECT 1.82 8.479 1.876 8.679 ;
 RECT 2.24 8.479 2.296 8.679 ;
 RECT 2.744 8.389 2.8 8.589 ;
 RECT 3.164 8.479 3.22 8.679 ;
 RECT 3.92 8.479 3.976 8.679 ;
 RECT 3.752 8.749 3.808 8.949 ;
 RECT 4.508 8.6785 4.564 8.8785 ;
 RECT 0.392 7.219 0.448 7.419 ;
 RECT 0.812 7.305 0.868 7.505 ;
 RECT 0.644 7.219 0.7 7.419 ;
 RECT 1.232 7.219 1.288 7.419 ;
 RECT 1.4 7.219 1.456 7.419 ;
 RECT 1.568 7.219 1.624 7.419 ;
 RECT 1.82 7.219 1.876 7.419 ;
 RECT 2.24 7.219 2.296 7.419 ;
 RECT 2.744 7.129 2.8 7.329 ;
 RECT 3.164 7.219 3.22 7.419 ;
 RECT 3.92 7.219 3.976 7.419 ;
 RECT 3.752 7.489 3.808 7.689 ;
 RECT 4.508 7.4185 4.564 7.6185 ;
 RECT 0.392 5.959 0.448 6.159 ;
 RECT 0.812 6.045 0.868 6.245 ;
 RECT 0.644 5.959 0.7 6.159 ;
 RECT 1.232 5.959 1.288 6.159 ;
 RECT 1.4 5.959 1.456 6.159 ;
 RECT 1.568 5.959 1.624 6.159 ;
 RECT 1.82 5.959 1.876 6.159 ;
 RECT 2.24 5.959 2.296 6.159 ;
 RECT 2.744 5.869 2.8 6.069 ;
 RECT 3.164 5.959 3.22 6.159 ;
 RECT 3.92 5.959 3.976 6.159 ;
 RECT 3.752 6.229 3.808 6.429 ;
 RECT 4.508 6.1585 4.564 6.3585 ;
 END
 END vss.gds444
 PIN vss.gds445
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.134 8.0595 10.194 8.2595 ;
 END
 END vss.gds445
 PIN vss.gds446
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.966 8.0595 10.026 8.2595 ;
 END
 END vss.gds446
 PIN vss.gds447
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.798 8.0595 9.858 8.2595 ;
 END
 END vss.gds447
 PIN vss.gds448
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.79 8.0595 8.85 8.2595 ;
 END
 END vss.gds448
 PIN vss.gds449
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.622 8.0595 8.682 8.2595 ;
 END
 END vss.gds449
 PIN vss.gds450
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.454 8.0595 8.514 8.2595 ;
 END
 END vss.gds450
 PIN vss.gds451
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 8.0595 9.69 8.2595 ;
 END
 END vss.gds451
 PIN vss.gds452
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.118 8.0595 8.178 8.2595 ;
 END
 END vss.gds452
 PIN vss.gds453
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 8.0595 8.346 8.2595 ;
 END
 END vss.gds453
 PIN vss.gds454
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.95 8.0595 8.01 8.2595 ;
 END
 END vss.gds454
 PIN vss.gds455
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.782 8.0595 7.842 8.2595 ;
 END
 END vss.gds455
 PIN vss.gds456
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.462 8.0595 9.522 8.2595 ;
 END
 END vss.gds456
 PIN vss.gds457
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.294 8.0595 9.354 8.2595 ;
 END
 END vss.gds457
 PIN vss.gds458
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.126 8.0595 9.186 8.2595 ;
 END
 END vss.gds458
 PIN vss.gds459
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.446 8.0595 7.506 8.2595 ;
 END
 END vss.gds459
 PIN vss.gds460
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 8.0595 9.018 8.2595 ;
 END
 END vss.gds460
 PIN vss.gds461
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 8.0595 7.674 8.2595 ;
 END
 END vss.gds461
 PIN vss.gds462
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 8.831 5.474 9.031 ;
 END
 END vss.gds462
 PIN vss.gds463
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 7.843 5.986 8.043 ;
 END
 END vss.gds463
 PIN vss.gds464
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 8.831 5.73 9.031 ;
 END
 END vss.gds464
 PIN vss.gds465
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.278 8.0595 7.338 8.2595 ;
 END
 END vss.gds465
 PIN vss.gds466
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.11 8.0595 7.17 8.2595 ;
 END
 END vss.gds466
 PIN vss.gds467
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 7.639 6.434 7.839 ;
 END
 END vss.gds467
 PIN vss.gds468
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 7.64 6.178 7.84 ;
 END
 END vss.gds468
 PIN vss.gds469
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 6.524 9.701 6.58 9.901 ;
 RECT 6.524 8.441 6.58 8.641 ;
 RECT 6.524 7.181 6.58 7.381 ;
 RECT 6.524 5.921 6.58 6.121 ;
 RECT 6.692 10.024 6.748 10.224 ;
 RECT 6.692 8.764 6.748 8.964 ;
 RECT 6.692 7.504 6.748 7.704 ;
 RECT 6.692 6.244 6.748 6.444 ;
 RECT 6.608 10.009 6.664 10.209 ;
 RECT 6.608 8.749 6.664 8.949 ;
 RECT 6.608 7.489 6.664 7.689 ;
 RECT 6.608 6.229 6.664 6.429 ;
 END
 END vss.gds469
 PIN vss.gds470
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 9.018 14.87 9.218 ;
 END
 END vss.gds470
 PIN vss.gds471
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 7.718 13.898 7.918 ;
 END
 END vss.gds471
 PIN vss.gds472
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 7.758 14.87 7.958 ;
 END
 END vss.gds472
 PIN vss.gds473
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 6.458 13.898 6.658 ;
 END
 END vss.gds473
 PIN vss.gds474
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 6.498 14.87 6.698 ;
 END
 END vss.gds474
 PIN vss.gds475
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.15 8.0595 12.21 8.2595 ;
 END
 END vss.gds475
 PIN vss.gds476
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.982 8.0595 12.042 8.2595 ;
 END
 END vss.gds476
 PIN vss.gds477
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.814 8.0595 11.874 8.2595 ;
 END
 END vss.gds477
 PIN vss.gds478
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 8.0595 13.658 8.2595 ;
 END
 END vss.gds478
 PIN vss.gds479
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 8.0595 11.706 8.2595 ;
 END
 END vss.gds479
 PIN vss.gds480
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.478 8.0595 11.538 8.2595 ;
 END
 END vss.gds480
 PIN vss.gds481
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.31 8.0595 11.37 8.2595 ;
 END
 END vss.gds481
 PIN vss.gds482
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.142 8.0595 11.202 8.2595 ;
 END
 END vss.gds482
 PIN vss.gds483
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.806 8.0595 10.866 8.2595 ;
 END
 END vss.gds483
 PIN vss.gds484
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.638 8.0595 10.698 8.2595 ;
 END
 END vss.gds484
 PIN vss.gds485
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.47 8.0595 10.53 8.2595 ;
 END
 END vss.gds485
 PIN vss.gds486
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 8.0595 11.034 8.2595 ;
 END
 END vss.gds486
 PIN vss.gds487
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 8.1 15.162 8.3 ;
 END
 END vss.gds487
 PIN vss.gds488
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 8.0595 10.362 8.2595 ;
 END
 END vss.gds488
 PIN vss.gds489
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 8.1 14.498 8.3 ;
 END
 END vss.gds489
 PIN vss.gds490
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 8.978 13.898 9.178 ;
 END
 END vss.gds490
 PIN vss.gds491
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.262 8.112 13.318 8.312 ;
 END
 END vss.gds491
 PIN vss.gds492
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 7.9635 12.818 8.1635 ;
 END
 END vss.gds492
 PIN vss.gds493
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 7.981 12.378 8.181 ;
 END
 END vss.gds493
 PIN vss.gds494
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 8.831 12.59 9.031 ;
 END
 END vss.gds494
 PIN vss.gds495
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 8.6535 13.058 8.8535 ;
 END
 END vss.gds495
 PIN vss.gds496
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 10.238 13.898 10.438 ;
 END
 END vss.gds496
 PIN vss.gds497
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 14 10.416 14.056 10.589 ;
 RECT 14.168 10.389 14.224 10.589 ;
 RECT 14 6.636 14.056 6.809 ;
 RECT 14.168 6.609 14.224 6.809 ;
 RECT 14 7.896 14.056 8.069 ;
 RECT 14.168 7.869 14.224 8.069 ;
 RECT 14 9.156 14.056 9.329 ;
 RECT 14.168 9.129 14.224 9.329 ;
 RECT 14.336 7.229 14.392 7.429 ;
 RECT 14.168 7.229 14.224 7.429 ;
 RECT 14.336 5.969 14.392 6.169 ;
 RECT 14.168 5.969 14.224 6.169 ;
 RECT 14.336 8.489 14.392 8.689 ;
 RECT 14.168 8.489 14.224 8.689 ;
 RECT 13.664 8.623 13.72 8.823 ;
 RECT 14.84 9.173 14.896 9.338 ;
 RECT 14.672 9.173 14.728 9.338 ;
 RECT 15.008 8.699 15.064 8.899 ;
 RECT 15.008 7.439 15.064 7.639 ;
 RECT 14.84 7.913 14.896 8.078 ;
 RECT 14.672 7.913 14.728 8.078 ;
 RECT 13.664 7.363 13.72 7.563 ;
 RECT 15.008 6.179 15.064 6.379 ;
 RECT 14.84 6.653 14.896 6.818 ;
 RECT 14.672 6.653 14.728 6.818 ;
 RECT 13.664 6.103 13.72 6.303 ;
 RECT 14.336 9.749 14.392 9.949 ;
 RECT 14.168 9.749 14.224 9.949 ;
 RECT 15.008 9.959 15.064 10.159 ;
 RECT 14.84 10.433 14.896 10.598 ;
 RECT 14.672 10.433 14.728 10.598 ;
 RECT 13.664 9.883 13.72 10.083 ;
 RECT 15.176 8.1395 15.232 8.3395 ;
 RECT 12.824 7.924 12.88 8.124 ;
 RECT 13.496 7.935 13.552 8.135 ;
 RECT 13.328 7.873 13.384 8.073 ;
 RECT 13.16 7.924 13.216 8.124 ;
 RECT 12.488 7.954 12.544 8.154 ;
 RECT 12.992 7.924 13.048 8.124 ;
 RECT 12.656 7.954 12.712 8.154 ;
 END
 END vss.gds497
 PIN vss.gds498
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.986 7.843 18.026 8.043 ;
 END
 END vss.gds498
 PIN vss.gds499
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.206 8.0595 19.266 8.2595 ;
 END
 END vss.gds499
 PIN vss.gds500
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.038 8.0595 19.098 8.2595 ;
 END
 END vss.gds500
 PIN vss.gds501
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.702 8.0595 18.762 8.2595 ;
 END
 END vss.gds501
 PIN vss.gds502
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 8.0595 20.274 8.2595 ;
 END
 END vss.gds502
 PIN vss.gds503
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.374 8.0595 19.434 8.2595 ;
 END
 END vss.gds503
 PIN vss.gds504
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 8.112 16.814 8.312 ;
 END
 END vss.gds504
 PIN vss.gds505
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 9.733 16.146 9.933 ;
 END
 END vss.gds505
 PIN vss.gds506
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 7.956 15.418 8.156 ;
 END
 END vss.gds506
 PIN vss.gds507
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 8.0595 19.602 8.2595 ;
 END
 END vss.gds507
 PIN vss.gds508
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 8.0595 18.93 8.2595 ;
 END
 END vss.gds508
 PIN vss.gds509
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 8.0185 16.994 8.2185 ;
 END
 END vss.gds509
 PIN vss.gds510
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 8.473 16.146 8.673 ;
 END
 END vss.gds510
 PIN vss.gds511
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 7.213 16.146 7.413 ;
 END
 END vss.gds511
 PIN vss.gds512
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 8.1 15.842 8.3 ;
 END
 END vss.gds512
 PIN vss.gds513
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.534 8.0595 18.594 8.2595 ;
 END
 END vss.gds513
 PIN vss.gds514
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 5.953 16.146 6.153 ;
 END
 END vss.gds514
 PIN vss.gds515
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.71 8.0595 19.77 8.2595 ;
 END
 END vss.gds515
 PIN vss.gds516
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.878 8.0595 19.938 8.2595 ;
 END
 END vss.gds516
 PIN vss.gds517
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 7.9635 17.834 8.1635 ;
 END
 END vss.gds517
 PIN vss.gds518
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.438 8.1155 17.494 8.3155 ;
 END
 END vss.gds518
 PIN vss.gds519
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.366 8.0595 18.426 8.2595 ;
 END
 END vss.gds519
 PIN vss.gds520
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.046 8.0595 20.106 8.2595 ;
 END
 END vss.gds520
 PIN vss.gds521
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 7.8665 16.49 8.0665 ;
 END
 END vss.gds521
 PIN vss.gds522
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 7.981 18.258 8.181 ;
 END
 END vss.gds522
 PIN vss.gds523
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 7.9635 17.314 8.1635 ;
 END
 END vss.gds523
 PIN vss.gds524
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 15.596 9.4 15.652 9.6 ;
 RECT 15.848 9.403 15.904 9.603 ;
 RECT 16.52 10.436 16.576 10.589 ;
 RECT 15.764 10.433 15.82 10.598 ;
 RECT 15.596 10.433 15.652 10.598 ;
 RECT 15.596 5.62 15.652 5.82 ;
 RECT 15.848 5.623 15.904 5.823 ;
 RECT 16.52 6.656 16.576 6.809 ;
 RECT 15.764 6.653 15.82 6.818 ;
 RECT 15.596 6.653 15.652 6.818 ;
 RECT 15.596 6.88 15.652 7.08 ;
 RECT 15.848 6.883 15.904 7.083 ;
 RECT 16.52 7.916 16.576 8.069 ;
 RECT 15.764 7.913 15.82 8.078 ;
 RECT 15.596 7.913 15.652 8.078 ;
 RECT 15.596 8.14 15.652 8.34 ;
 RECT 15.848 8.143 15.904 8.343 ;
 RECT 16.52 9.176 16.576 9.329 ;
 RECT 16.352 8.7995 16.408 8.9995 ;
 RECT 16.856 8.5475 16.912 8.7475 ;
 RECT 15.764 9.173 15.82 9.338 ;
 RECT 15.596 9.173 15.652 9.338 ;
 RECT 15.428 8.699 15.484 8.899 ;
 RECT 15.428 7.439 15.484 7.639 ;
 RECT 16.856 7.2875 16.912 7.4875 ;
 RECT 16.352 7.5395 16.408 7.7395 ;
 RECT 15.428 6.179 15.484 6.379 ;
 RECT 16.352 6.2795 16.408 6.4795 ;
 RECT 16.856 6.0275 16.912 6.2275 ;
 RECT 15.428 9.959 15.484 10.159 ;
 RECT 16.856 9.8075 16.912 10.0075 ;
 RECT 16.352 10.0595 16.408 10.2595 ;
 RECT 17.864 7.954 17.92 8.154 ;
 RECT 17.696 7.9615 17.752 8.1615 ;
 RECT 17.528 7.954 17.584 8.154 ;
 RECT 17.36 7.954 17.416 8.154 ;
 RECT 17.192 7.954 17.248 8.154 ;
 RECT 17.024 8.069 17.08 8.269 ;
 RECT 18.032 7.954 18.088 8.154 ;
 END
 END vss.gds524
 PIN vss.gds525
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.17 8.0595 25.23 8.2595 ;
 END
 END vss.gds525
 PIN vss.gds526
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.002 8.0595 25.062 8.2595 ;
 END
 END vss.gds526
 PIN vss.gds527
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.834 8.0595 24.894 8.2595 ;
 END
 END vss.gds527
 PIN vss.gds528
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.498 8.0595 24.558 8.2595 ;
 END
 END vss.gds528
 PIN vss.gds529
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.33 8.0595 24.39 8.2595 ;
 END
 END vss.gds529
 PIN vss.gds530
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.162 8.0595 24.222 8.2595 ;
 END
 END vss.gds530
 PIN vss.gds531
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.406 8.0595 23.466 8.2595 ;
 END
 END vss.gds531
 PIN vss.gds532
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.238 8.0595 23.298 8.2595 ;
 END
 END vss.gds532
 PIN vss.gds533
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.07 8.0595 23.13 8.2595 ;
 END
 END vss.gds533
 PIN vss.gds534
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.734 8.0595 22.794 8.2595 ;
 END
 END vss.gds534
 PIN vss.gds535
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.566 8.0595 22.626 8.2595 ;
 END
 END vss.gds535
 PIN vss.gds536
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.398 8.0595 22.458 8.2595 ;
 END
 END vss.gds536
 PIN vss.gds537
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.062 8.0595 22.122 8.2595 ;
 END
 END vss.gds537
 PIN vss.gds538
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.894 8.0595 21.954 8.2595 ;
 END
 END vss.gds538
 PIN vss.gds539
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.726 8.0595 21.786 8.2595 ;
 END
 END vss.gds539
 PIN vss.gds540
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.39 8.0595 21.45 8.2595 ;
 END
 END vss.gds540
 PIN vss.gds541
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.222 8.0595 21.282 8.2595 ;
 END
 END vss.gds541
 PIN vss.gds542
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.054 8.0595 21.114 8.2595 ;
 END
 END vss.gds542
 PIN vss.gds543
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.718 8.0595 20.778 8.2595 ;
 END
 END vss.gds543
 PIN vss.gds544
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.55 8.0595 20.61 8.2595 ;
 END
 END vss.gds544
 PIN vss.gds545
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.382 8.0595 20.442 8.2595 ;
 END
 END vss.gds545
 PIN vss.gds546
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 8.0595 24.726 8.2595 ;
 END
 END vss.gds546
 PIN vss.gds547
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 8.0595 22.962 8.2595 ;
 END
 END vss.gds547
 PIN vss.gds548
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 8.0595 22.29 8.2595 ;
 END
 END vss.gds548
 PIN vss.gds549
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 8.0595 21.618 8.2595 ;
 END
 END vss.gds549
 PIN vss.gds550
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 8.0595 20.946 8.2595 ;
 END
 END vss.gds550
 PIN vss.gds551
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 8.0595 23.634 8.2595 ;
 END
 END vss.gds551
 PIN vss.gds552
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 23.912 8.636 23.968 8.836 ;
 RECT 23.912 7.376 23.968 7.576 ;
 RECT 23.912 6.116 23.968 6.316 ;
 RECT 23.912 9.896 23.968 10.096 ;
 RECT 23.744 8.006 23.8 8.206 ;
 END
 END vss.gds552
 PIN vss.gds553
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.202 8.0595 29.262 8.2595 ;
 END
 END vss.gds553
 PIN vss.gds554
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.034 8.0595 29.094 8.2595 ;
 END
 END vss.gds554
 PIN vss.gds555
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.866 8.0595 28.926 8.2595 ;
 END
 END vss.gds555
 PIN vss.gds556
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.53 8.0595 28.59 8.2595 ;
 END
 END vss.gds556
 PIN vss.gds557
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.362 8.0595 28.422 8.2595 ;
 END
 END vss.gds557
 PIN vss.gds558
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.194 8.0595 28.254 8.2595 ;
 END
 END vss.gds558
 PIN vss.gds559
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.858 8.0595 27.918 8.2595 ;
 END
 END vss.gds559
 PIN vss.gds560
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.69 8.0595 27.75 8.2595 ;
 END
 END vss.gds560
 PIN vss.gds561
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.522 8.0595 27.582 8.2595 ;
 END
 END vss.gds561
 PIN vss.gds562
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.186 8.0595 27.246 8.2595 ;
 END
 END vss.gds562
 PIN vss.gds563
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.018 8.0595 27.078 8.2595 ;
 END
 END vss.gds563
 PIN vss.gds564
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.85 8.0595 26.91 8.2595 ;
 END
 END vss.gds564
 PIN vss.gds565
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.514 8.0595 26.574 8.2595 ;
 END
 END vss.gds565
 PIN vss.gds566
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.346 8.0595 26.406 8.2595 ;
 END
 END vss.gds566
 PIN vss.gds567
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.178 8.0595 26.238 8.2595 ;
 END
 END vss.gds567
 PIN vss.gds568
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.842 8.0595 25.902 8.2595 ;
 END
 END vss.gds568
 PIN vss.gds569
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.674 8.0595 25.734 8.2595 ;
 END
 END vss.gds569
 PIN vss.gds570
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.506 8.0595 25.566 8.2595 ;
 END
 END vss.gds570
 PIN vss.gds571
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 8.6535 30.11 8.8535 ;
 END
 END vss.gds571
 PIN vss.gds572
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 7.981 29.43 8.181 ;
 END
 END vss.gds572
 PIN vss.gds573
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 8.0595 28.758 8.2595 ;
 END
 END vss.gds573
 PIN vss.gds574
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 8.0595 28.086 8.2595 ;
 END
 END vss.gds574
 PIN vss.gds575
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 8.0595 27.414 8.2595 ;
 END
 END vss.gds575
 PIN vss.gds576
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 8.0595 26.742 8.2595 ;
 END
 END vss.gds576
 PIN vss.gds577
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 8.0595 26.07 8.2595 ;
 END
 END vss.gds577
 PIN vss.gds578
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 8.0595 25.398 8.2595 ;
 END
 END vss.gds578
 PIN vss.gds579
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 7.9635 29.87 8.1635 ;
 END
 END vss.gds579
 PIN vss.gds580
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 8.831 29.642 9.031 ;
 END
 END vss.gds580
 PIN vss.gds581
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.876 7.924 29.932 8.124 ;
 RECT 29.54 7.954 29.596 8.154 ;
 RECT 30.212 7.924 30.268 8.124 ;
 RECT 30.044 7.924 30.1 8.124 ;
 RECT 29.708 7.954 29.764 8.154 ;
 END
 END vss.gds581
 PIN vss.gds582
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 9.018 31.922 9.218 ;
 END
 END vss.gds582
 PIN vss.gds583
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 8.978 30.95 9.178 ;
 END
 END vss.gds583
 PIN vss.gds584
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.038 7.843 35.078 8.043 ;
 END
 END vss.gds584
 PIN vss.gds585
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 7.718 30.95 7.918 ;
 END
 END vss.gds585
 PIN vss.gds586
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 7.758 31.922 7.958 ;
 END
 END vss.gds586
 PIN vss.gds587
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 6.458 30.95 6.658 ;
 END
 END vss.gds587
 PIN vss.gds588
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 6.498 31.922 6.698 ;
 END
 END vss.gds588
 PIN vss.gds589
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.314 8.112 30.37 8.312 ;
 END
 END vss.gds589
 PIN vss.gds590
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 10.238 30.95 10.438 ;
 END
 END vss.gds590
 PIN vss.gds591
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 8.1 32.894 8.3 ;
 END
 END vss.gds591
 PIN vss.gds592
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 8.1 32.214 8.3 ;
 END
 END vss.gds592
 PIN vss.gds593
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 7.956 32.47 8.156 ;
 END
 END vss.gds593
 PIN vss.gds594
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 8.0595 30.71 8.2595 ;
 END
 END vss.gds594
 PIN vss.gds595
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 7.8665 33.542 8.0665 ;
 END
 END vss.gds595
 PIN vss.gds596
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 9.733 33.198 9.933 ;
 END
 END vss.gds596
 PIN vss.gds597
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 8.473 33.198 8.673 ;
 END
 END vss.gds597
 PIN vss.gds598
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 7.213 33.198 7.413 ;
 END
 END vss.gds598
 PIN vss.gds599
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 8.1 31.55 8.3 ;
 END
 END vss.gds599
 PIN vss.gds600
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 5.953 33.198 6.153 ;
 END
 END vss.gds600
 PIN vss.gds601
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 8.112 33.866 8.312 ;
 END
 END vss.gds601
 PIN vss.gds602
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 7.9635 34.886 8.1635 ;
 END
 END vss.gds602
 PIN vss.gds603
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.49 8.1155 34.546 8.3155 ;
 END
 END vss.gds603
 PIN vss.gds604
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 8.0185 34.046 8.2185 ;
 END
 END vss.gds604
 PIN vss.gds605
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 7.9635 34.366 8.1635 ;
 END
 END vss.gds605
 PIN vss.gds606
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 32.648 9.4 32.704 9.6 ;
 RECT 32.9 9.403 32.956 9.603 ;
 RECT 33.572 10.436 33.628 10.589 ;
 RECT 31.052 10.416 31.108 10.589 ;
 RECT 31.22 10.389 31.276 10.589 ;
 RECT 32.816 10.433 32.872 10.598 ;
 RECT 32.648 10.433 32.704 10.598 ;
 RECT 31.892 10.433 31.948 10.598 ;
 RECT 31.724 10.433 31.78 10.598 ;
 RECT 32.648 5.62 32.704 5.82 ;
 RECT 32.9 5.623 32.956 5.823 ;
 RECT 33.572 6.656 33.628 6.809 ;
 RECT 31.052 6.636 31.108 6.809 ;
 RECT 31.22 6.609 31.276 6.809 ;
 RECT 32.816 6.653 32.872 6.818 ;
 RECT 32.648 6.653 32.704 6.818 ;
 RECT 31.892 6.653 31.948 6.818 ;
 RECT 31.724 6.653 31.78 6.818 ;
 RECT 33.572 7.916 33.628 8.069 ;
 RECT 31.052 7.896 31.108 8.069 ;
 RECT 31.22 7.869 31.276 8.069 ;
 RECT 32.816 7.913 32.872 8.078 ;
 RECT 32.648 7.913 32.704 8.078 ;
 RECT 31.892 7.913 31.948 8.078 ;
 RECT 31.724 7.913 31.78 8.078 ;
 RECT 33.572 9.176 33.628 9.329 ;
 RECT 31.052 9.156 31.108 9.329 ;
 RECT 31.22 9.129 31.276 9.329 ;
 RECT 32.816 9.173 32.872 9.338 ;
 RECT 32.648 9.173 32.704 9.338 ;
 RECT 31.892 9.173 31.948 9.338 ;
 RECT 31.724 9.173 31.78 9.338 ;
 RECT 32.648 6.88 32.704 7.08 ;
 RECT 32.9 6.883 32.956 7.083 ;
 RECT 32.648 8.14 32.704 8.34 ;
 RECT 32.9 8.143 32.956 8.343 ;
 RECT 31.388 7.229 31.444 7.429 ;
 RECT 31.22 7.229 31.276 7.429 ;
 RECT 31.388 9.749 31.444 9.949 ;
 RECT 31.22 9.749 31.276 9.949 ;
 RECT 30.716 9.883 30.772 10.083 ;
 RECT 32.06 9.959 32.116 10.159 ;
 RECT 32.48 9.959 32.536 10.159 ;
 RECT 32.06 8.699 32.116 8.899 ;
 RECT 32.48 8.699 32.536 8.899 ;
 RECT 31.388 8.489 31.444 8.689 ;
 RECT 31.22 8.489 31.276 8.689 ;
 RECT 30.716 8.623 30.772 8.823 ;
 RECT 30.716 7.363 30.772 7.563 ;
 RECT 33.404 7.5395 33.46 7.7395 ;
 RECT 33.908 7.2875 33.964 7.4875 ;
 RECT 33.908 6.0275 33.964 6.2275 ;
 RECT 33.404 6.2795 33.46 6.4795 ;
 RECT 32.06 6.179 32.116 6.379 ;
 RECT 32.48 6.179 32.536 6.379 ;
 RECT 31.388 5.969 31.444 6.169 ;
 RECT 31.22 5.969 31.276 6.169 ;
 RECT 30.716 6.103 30.772 6.303 ;
 RECT 32.06 7.439 32.116 7.639 ;
 RECT 32.48 7.439 32.536 7.639 ;
 RECT 33.404 8.7995 33.46 8.9995 ;
 RECT 33.908 8.5475 33.964 8.7475 ;
 RECT 30.548 7.935 30.604 8.135 ;
 RECT 33.908 9.8075 33.964 10.0075 ;
 RECT 33.404 10.0595 33.46 10.2595 ;
 RECT 30.38 7.873 30.436 8.073 ;
 RECT 32.228 8.1395 32.284 8.3395 ;
 RECT 34.916 7.954 34.972 8.154 ;
 RECT 34.748 7.9615 34.804 8.1615 ;
 RECT 34.58 7.954 34.636 8.154 ;
 RECT 34.412 7.954 34.468 8.154 ;
 RECT 34.244 7.954 34.3 8.154 ;
 RECT 35.084 7.954 35.14 8.154 ;
 RECT 34.076 8.069 34.132 8.269 ;
 END
 END vss.gds606
 PIN vss.gds607
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.122 8.0595 40.182 8.2595 ;
 END
 END vss.gds607
 PIN vss.gds608
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.586 8.0595 35.646 8.2595 ;
 END
 END vss.gds608
 PIN vss.gds609
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.754 8.0595 35.814 8.2595 ;
 END
 END vss.gds609
 PIN vss.gds610
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.09 8.0595 36.15 8.2595 ;
 END
 END vss.gds610
 PIN vss.gds611
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.258 8.0595 36.318 8.2595 ;
 END
 END vss.gds611
 PIN vss.gds612
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.426 8.0595 36.486 8.2595 ;
 END
 END vss.gds612
 PIN vss.gds613
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.762 8.0595 36.822 8.2595 ;
 END
 END vss.gds613
 PIN vss.gds614
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.93 8.0595 36.99 8.2595 ;
 END
 END vss.gds614
 PIN vss.gds615
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.098 8.0595 37.158 8.2595 ;
 END
 END vss.gds615
 PIN vss.gds616
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.434 8.0595 37.494 8.2595 ;
 END
 END vss.gds616
 PIN vss.gds617
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.602 8.0595 37.662 8.2595 ;
 END
 END vss.gds617
 PIN vss.gds618
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.77 8.0595 37.83 8.2595 ;
 END
 END vss.gds618
 PIN vss.gds619
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.106 8.0595 38.166 8.2595 ;
 END
 END vss.gds619
 PIN vss.gds620
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.274 8.0595 38.334 8.2595 ;
 END
 END vss.gds620
 PIN vss.gds621
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.442 8.0595 38.502 8.2595 ;
 END
 END vss.gds621
 PIN vss.gds622
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.778 8.0595 38.838 8.2595 ;
 END
 END vss.gds622
 PIN vss.gds623
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.946 8.0595 39.006 8.2595 ;
 END
 END vss.gds623
 PIN vss.gds624
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 8.0595 37.998 8.2595 ;
 END
 END vss.gds624
 PIN vss.gds625
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 8.0595 37.326 8.2595 ;
 END
 END vss.gds625
 PIN vss.gds626
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 8.0595 38.67 8.2595 ;
 END
 END vss.gds626
 PIN vss.gds627
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.45 8.0595 39.51 8.2595 ;
 END
 END vss.gds627
 PIN vss.gds628
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 8.0595 36.654 8.2595 ;
 END
 END vss.gds628
 PIN vss.gds629
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.618 8.0595 39.678 8.2595 ;
 END
 END vss.gds629
 PIN vss.gds630
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.786 8.0595 39.846 8.2595 ;
 END
 END vss.gds630
 PIN vss.gds631
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 8.0595 39.342 8.2595 ;
 END
 END vss.gds631
 PIN vss.gds632
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.114 8.0595 39.174 8.2595 ;
 END
 END vss.gds632
 PIN vss.gds633
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 8.0595 40.014 8.2595 ;
 END
 END vss.gds633
 PIN vss.gds634
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.418 8.0595 35.478 8.2595 ;
 END
 END vss.gds634
 PIN vss.gds635
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 7.981 35.31 8.181 ;
 END
 END vss.gds635
 PIN vss.gds636
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 8.0595 35.982 8.2595 ;
 END
 END vss.gds636
 PIN vss.gds637
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.91 8.0595 44.97 8.2595 ;
 END
 END vss.gds637
 PIN vss.gds638
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.742 8.0595 44.802 8.2595 ;
 END
 END vss.gds638
 PIN vss.gds639
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.574 8.0595 44.634 8.2595 ;
 END
 END vss.gds639
 PIN vss.gds640
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.238 8.0595 44.298 8.2595 ;
 END
 END vss.gds640
 PIN vss.gds641
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.07 8.0595 44.13 8.2595 ;
 END
 END vss.gds641
 PIN vss.gds642
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.902 8.0595 43.962 8.2595 ;
 END
 END vss.gds642
 PIN vss.gds643
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.566 8.0595 43.626 8.2595 ;
 END
 END vss.gds643
 PIN vss.gds644
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.398 8.0595 43.458 8.2595 ;
 END
 END vss.gds644
 PIN vss.gds645
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.23 8.0595 43.29 8.2595 ;
 END
 END vss.gds645
 PIN vss.gds646
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.894 8.0595 42.954 8.2595 ;
 END
 END vss.gds646
 PIN vss.gds647
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.726 8.0595 42.786 8.2595 ;
 END
 END vss.gds647
 PIN vss.gds648
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.558 8.0595 42.618 8.2595 ;
 END
 END vss.gds648
 PIN vss.gds649
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.222 8.0595 42.282 8.2595 ;
 END
 END vss.gds649
 PIN vss.gds650
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.054 8.0595 42.114 8.2595 ;
 END
 END vss.gds650
 PIN vss.gds651
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.886 8.0595 41.946 8.2595 ;
 END
 END vss.gds651
 PIN vss.gds652
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.55 8.0595 41.61 8.2595 ;
 END
 END vss.gds652
 PIN vss.gds653
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.382 8.0595 41.442 8.2595 ;
 END
 END vss.gds653
 PIN vss.gds654
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.214 8.0595 41.274 8.2595 ;
 END
 END vss.gds654
 PIN vss.gds655
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.29 8.0595 40.35 8.2595 ;
 END
 END vss.gds655
 PIN vss.gds656
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.458 8.0595 40.518 8.2595 ;
 END
 END vss.gds656
 PIN vss.gds657
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 8.0595 45.138 8.2595 ;
 END
 END vss.gds657
 PIN vss.gds658
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 8.0595 44.466 8.2595 ;
 END
 END vss.gds658
 PIN vss.gds659
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 8.0595 43.794 8.2595 ;
 END
 END vss.gds659
 PIN vss.gds660
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 8.0595 43.122 8.2595 ;
 END
 END vss.gds660
 PIN vss.gds661
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 8.0595 42.45 8.2595 ;
 END
 END vss.gds661
 PIN vss.gds662
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 8.0595 41.778 8.2595 ;
 END
 END vss.gds662
 PIN vss.gds663
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 8.0595 40.686 8.2595 ;
 END
 END vss.gds663
 PIN vss.gds664
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 40.964 7.376 41.02 7.576 ;
 RECT 40.964 8.636 41.02 8.836 ;
 RECT 40.964 6.116 41.02 6.316 ;
 RECT 40.964 9.896 41.02 10.096 ;
 RECT 40.796 8.006 40.852 8.206 ;
 END
 END vss.gds664
 PIN vss.gds665
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 10.238 48.002 10.438 ;
 END
 END vss.gds665
 PIN vss.gds666
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 9.018 48.974 9.218 ;
 END
 END vss.gds666
 PIN vss.gds667
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 7.758 48.974 7.958 ;
 END
 END vss.gds667
 PIN vss.gds668
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 6.458 48.002 6.658 ;
 END
 END vss.gds668
 PIN vss.gds669
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 6.498 48.974 6.698 ;
 END
 END vss.gds669
 PIN vss.gds670
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 8.978 48.002 9.178 ;
 END
 END vss.gds670
 PIN vss.gds671
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.366 8.112 47.422 8.312 ;
 END
 END vss.gds671
 PIN vss.gds672
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.254 8.0595 46.314 8.2595 ;
 END
 END vss.gds672
 PIN vss.gds673
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.086 8.0595 46.146 8.2595 ;
 END
 END vss.gds673
 PIN vss.gds674
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.918 8.0595 45.978 8.2595 ;
 END
 END vss.gds674
 PIN vss.gds675
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.582 8.0595 45.642 8.2595 ;
 END
 END vss.gds675
 PIN vss.gds676
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.414 8.0595 45.474 8.2595 ;
 END
 END vss.gds676
 PIN vss.gds677
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.246 8.0595 45.306 8.2595 ;
 END
 END vss.gds677
 PIN vss.gds678
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 8.0595 45.81 8.2595 ;
 END
 END vss.gds678
 PIN vss.gds679
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 7.981 46.482 8.181 ;
 END
 END vss.gds679
 PIN vss.gds680
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 8.6535 47.162 8.8535 ;
 END
 END vss.gds680
 PIN vss.gds681
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 7.9635 46.922 8.1635 ;
 END
 END vss.gds681
 PIN vss.gds682
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 8.831 46.694 9.031 ;
 END
 END vss.gds682
 PIN vss.gds683
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 8.0595 47.762 8.2595 ;
 END
 END vss.gds683
 PIN vss.gds684
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 8.1 49.266 8.3 ;
 END
 END vss.gds684
 PIN vss.gds685
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 8.473 50.25 8.673 ;
 END
 END vss.gds685
 PIN vss.gds686
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 7.213 50.25 7.413 ;
 END
 END vss.gds686
 PIN vss.gds687
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 9.733 50.25 9.933 ;
 END
 END vss.gds687
 PIN vss.gds688
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 5.953 50.25 6.153 ;
 END
 END vss.gds688
 PIN vss.gds689
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 8.1 48.602 8.3 ;
 END
 END vss.gds689
 PIN vss.gds690
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 8.1 49.946 8.3 ;
 END
 END vss.gds690
 PIN vss.gds691
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 7.718 48.002 7.918 ;
 END
 END vss.gds691
 PIN vss.gds692
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 7.956 49.522 8.156 ;
 END
 END vss.gds692
 PIN vss.gds693
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 49.7 9.4 49.756 9.6 ;
 RECT 49.952 9.403 50.008 9.603 ;
 RECT 48.104 10.416 48.16 10.589 ;
 RECT 48.272 10.389 48.328 10.589 ;
 RECT 49.868 10.433 49.924 10.598 ;
 RECT 49.7 10.433 49.756 10.598 ;
 RECT 48.944 10.433 49 10.598 ;
 RECT 48.776 10.433 48.832 10.598 ;
 RECT 48.44 9.749 48.496 9.949 ;
 RECT 48.272 9.749 48.328 9.949 ;
 RECT 47.768 9.883 47.824 10.083 ;
 RECT 49.7 8.14 49.756 8.34 ;
 RECT 49.952 8.143 50.008 8.343 ;
 RECT 48.104 6.636 48.16 6.809 ;
 RECT 48.272 6.609 48.328 6.809 ;
 RECT 49.868 6.653 49.924 6.818 ;
 RECT 49.7 6.653 49.756 6.818 ;
 RECT 48.944 6.653 49 6.818 ;
 RECT 48.776 6.653 48.832 6.818 ;
 RECT 48.104 7.896 48.16 8.069 ;
 RECT 48.272 7.869 48.328 8.069 ;
 RECT 49.868 7.913 49.924 8.078 ;
 RECT 49.7 7.913 49.756 8.078 ;
 RECT 48.944 7.913 49 8.078 ;
 RECT 48.776 7.913 48.832 8.078 ;
 RECT 48.104 9.156 48.16 9.329 ;
 RECT 48.272 9.129 48.328 9.329 ;
 RECT 49.868 9.173 49.924 9.338 ;
 RECT 49.7 9.173 49.756 9.338 ;
 RECT 48.944 9.173 49 9.338 ;
 RECT 48.776 9.173 48.832 9.338 ;
 RECT 49.7 5.62 49.756 5.82 ;
 RECT 49.952 5.623 50.008 5.823 ;
 RECT 49.7 6.88 49.756 7.08 ;
 RECT 49.952 6.883 50.008 7.083 ;
 RECT 49.112 9.959 49.168 10.159 ;
 RECT 49.532 9.959 49.588 10.159 ;
 RECT 48.44 7.229 48.496 7.429 ;
 RECT 48.272 7.229 48.328 7.429 ;
 RECT 49.112 7.439 49.168 7.639 ;
 RECT 49.532 7.439 49.588 7.639 ;
 RECT 49.112 8.699 49.168 8.899 ;
 RECT 49.532 8.699 49.588 8.899 ;
 RECT 48.44 8.489 48.496 8.689 ;
 RECT 48.272 8.489 48.328 8.689 ;
 RECT 47.768 8.623 47.824 8.823 ;
 RECT 47.768 7.363 47.824 7.563 ;
 RECT 49.112 6.179 49.168 6.379 ;
 RECT 49.532 6.179 49.588 6.379 ;
 RECT 48.44 5.969 48.496 6.169 ;
 RECT 48.272 5.969 48.328 6.169 ;
 RECT 47.768 6.103 47.824 6.303 ;
 RECT 47.6 7.935 47.656 8.135 ;
 RECT 47.432 7.873 47.488 8.073 ;
 RECT 47.264 7.924 47.32 8.124 ;
 RECT 46.928 7.924 46.984 8.124 ;
 RECT 46.592 7.954 46.648 8.154 ;
 RECT 47.096 7.924 47.152 8.124 ;
 RECT 49.28 8.1395 49.336 8.3395 ;
 RECT 46.76 7.954 46.816 8.154 ;
 END
 END vss.gds693
 PIN vss.gds694
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.09 7.843 52.13 8.043 ;
 END
 END vss.gds694
 PIN vss.gds695
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.638 8.0595 52.698 8.2595 ;
 END
 END vss.gds695
 PIN vss.gds696
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.806 8.0595 52.866 8.2595 ;
 END
 END vss.gds696
 PIN vss.gds697
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.142 8.0595 53.202 8.2595 ;
 END
 END vss.gds697
 PIN vss.gds698
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.31 8.0595 53.37 8.2595 ;
 END
 END vss.gds698
 PIN vss.gds699
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.478 8.0595 53.538 8.2595 ;
 END
 END vss.gds699
 PIN vss.gds700
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.814 8.0595 53.874 8.2595 ;
 END
 END vss.gds700
 PIN vss.gds701
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.982 8.0595 54.042 8.2595 ;
 END
 END vss.gds701
 PIN vss.gds702
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.15 8.0595 54.21 8.2595 ;
 END
 END vss.gds702
 PIN vss.gds703
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.486 8.0595 54.546 8.2595 ;
 END
 END vss.gds703
 PIN vss.gds704
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.654 8.0595 54.714 8.2595 ;
 END
 END vss.gds704
 PIN vss.gds705
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.822 8.0595 54.882 8.2595 ;
 END
 END vss.gds705
 PIN vss.gds706
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.158 8.0595 55.218 8.2595 ;
 END
 END vss.gds706
 PIN vss.gds707
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 8.0595 54.378 8.2595 ;
 END
 END vss.gds707
 PIN vss.gds708
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 8.0595 55.05 8.2595 ;
 END
 END vss.gds708
 PIN vss.gds709
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 8.0595 53.706 8.2595 ;
 END
 END vss.gds709
 PIN vss.gds710
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 7.9635 51.418 8.1635 ;
 END
 END vss.gds710
 PIN vss.gds711
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 8.112 50.918 8.312 ;
 END
 END vss.gds711
 PIN vss.gds712
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 8.0595 53.034 8.2595 ;
 END
 END vss.gds712
 PIN vss.gds713
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 7.9635 51.938 8.1635 ;
 END
 END vss.gds713
 PIN vss.gds714
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 7.8665 50.594 8.0665 ;
 END
 END vss.gds714
 PIN vss.gds715
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.47 8.0595 52.53 8.2595 ;
 END
 END vss.gds715
 PIN vss.gds716
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.542 8.1155 51.598 8.3155 ;
 END
 END vss.gds716
 PIN vss.gds717
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 7.981 52.362 8.181 ;
 END
 END vss.gds717
 PIN vss.gds718
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 8.0185 51.098 8.2185 ;
 END
 END vss.gds718
 PIN vss.gds719
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 50.624 10.436 50.68 10.589 ;
 RECT 50.624 6.656 50.68 6.809 ;
 RECT 50.624 7.916 50.68 8.069 ;
 RECT 50.624 9.176 50.68 9.329 ;
 RECT 50.456 7.5395 50.512 7.7395 ;
 RECT 50.96 7.2875 51.016 7.4875 ;
 RECT 50.96 8.5475 51.016 8.7475 ;
 RECT 50.456 8.7995 50.512 8.9995 ;
 RECT 50.96 6.0275 51.016 6.2275 ;
 RECT 50.456 6.2795 50.512 6.4795 ;
 RECT 50.96 9.8075 51.016 10.0075 ;
 RECT 50.456 10.0595 50.512 10.2595 ;
 RECT 51.968 7.954 52.024 8.154 ;
 RECT 51.8 7.9615 51.856 8.1615 ;
 RECT 51.632 7.954 51.688 8.154 ;
 RECT 51.464 7.954 51.52 8.154 ;
 RECT 51.296 7.954 51.352 8.154 ;
 RECT 52.136 7.954 52.192 8.154 ;
 RECT 51.128 8.069 51.184 8.269 ;
 END
 END vss.gds719
 PIN vss.gds720
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.946 8.0595 60.006 8.2595 ;
 END
 END vss.gds720
 PIN vss.gds721
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.778 8.0595 59.838 8.2595 ;
 END
 END vss.gds721
 PIN vss.gds722
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.61 8.0595 59.67 8.2595 ;
 END
 END vss.gds722
 PIN vss.gds723
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.274 8.0595 59.334 8.2595 ;
 END
 END vss.gds723
 PIN vss.gds724
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.106 8.0595 59.166 8.2595 ;
 END
 END vss.gds724
 PIN vss.gds725
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.938 8.0595 58.998 8.2595 ;
 END
 END vss.gds725
 PIN vss.gds726
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.602 8.0595 58.662 8.2595 ;
 END
 END vss.gds726
 PIN vss.gds727
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.434 8.0595 58.494 8.2595 ;
 END
 END vss.gds727
 PIN vss.gds728
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.266 8.0595 58.326 8.2595 ;
 END
 END vss.gds728
 PIN vss.gds729
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.326 8.0595 55.386 8.2595 ;
 END
 END vss.gds729
 PIN vss.gds730
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.494 8.0595 55.554 8.2595 ;
 END
 END vss.gds730
 PIN vss.gds731
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.83 8.0595 55.89 8.2595 ;
 END
 END vss.gds731
 PIN vss.gds732
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.998 8.0595 56.058 8.2595 ;
 END
 END vss.gds732
 PIN vss.gds733
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.166 8.0595 56.226 8.2595 ;
 END
 END vss.gds733
 PIN vss.gds734
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 8.0595 60.174 8.2595 ;
 END
 END vss.gds734
 PIN vss.gds735
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 8.0595 59.502 8.2595 ;
 END
 END vss.gds735
 PIN vss.gds736
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 8.0595 58.83 8.2595 ;
 END
 END vss.gds736
 PIN vss.gds737
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 8.0595 55.722 8.2595 ;
 END
 END vss.gds737
 PIN vss.gds738
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 8.0595 56.394 8.2595 ;
 END
 END vss.gds738
 PIN vss.gds739
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.502 8.0595 56.562 8.2595 ;
 END
 END vss.gds739
 PIN vss.gds740
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.67 8.0595 56.73 8.2595 ;
 END
 END vss.gds740
 PIN vss.gds741
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.838 8.0595 56.898 8.2595 ;
 END
 END vss.gds741
 PIN vss.gds742
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.342 8.0595 57.402 8.2595 ;
 END
 END vss.gds742
 PIN vss.gds743
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.51 8.0595 57.57 8.2595 ;
 END
 END vss.gds743
 PIN vss.gds744
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 8.0595 57.738 8.2595 ;
 END
 END vss.gds744
 PIN vss.gds745
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 8.0595 57.066 8.2595 ;
 END
 END vss.gds745
 PIN vss.gds746
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.174 8.0595 57.234 8.2595 ;
 END
 END vss.gds746
 PIN vss.gds747
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 58.016 7.376 58.072 7.576 ;
 RECT 58.016 8.636 58.072 8.836 ;
 RECT 58.016 6.116 58.072 6.316 ;
 RECT 58.016 9.896 58.072 10.096 ;
 RECT 57.848 8.006 57.904 8.206 ;
 END
 END vss.gds747
 PIN vss.gds748
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 10.238 65.054 10.438 ;
 END
 END vss.gds748
 PIN vss.gds749
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 7.718 65.054 7.918 ;
 END
 END vss.gds749
 PIN vss.gds750
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 8.978 65.054 9.178 ;
 END
 END vss.gds750
 PIN vss.gds751
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.418 8.112 64.474 8.312 ;
 END
 END vss.gds751
 PIN vss.gds752
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.306 8.0595 63.366 8.2595 ;
 END
 END vss.gds752
 PIN vss.gds753
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.138 8.0595 63.198 8.2595 ;
 END
 END vss.gds753
 PIN vss.gds754
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.97 8.0595 63.03 8.2595 ;
 END
 END vss.gds754
 PIN vss.gds755
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.634 8.0595 62.694 8.2595 ;
 END
 END vss.gds755
 PIN vss.gds756
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.466 8.0595 62.526 8.2595 ;
 END
 END vss.gds756
 PIN vss.gds757
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.298 8.0595 62.358 8.2595 ;
 END
 END vss.gds757
 PIN vss.gds758
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.962 8.0595 62.022 8.2595 ;
 END
 END vss.gds758
 PIN vss.gds759
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.794 8.0595 61.854 8.2595 ;
 END
 END vss.gds759
 PIN vss.gds760
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.626 8.0595 61.686 8.2595 ;
 END
 END vss.gds760
 PIN vss.gds761
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.29 8.0595 61.35 8.2595 ;
 END
 END vss.gds761
 PIN vss.gds762
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.122 8.0595 61.182 8.2595 ;
 END
 END vss.gds762
 PIN vss.gds763
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.954 8.0595 61.014 8.2595 ;
 END
 END vss.gds763
 PIN vss.gds764
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.618 8.0595 60.678 8.2595 ;
 END
 END vss.gds764
 PIN vss.gds765
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.45 8.0595 60.51 8.2595 ;
 END
 END vss.gds765
 PIN vss.gds766
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.282 8.0595 60.342 8.2595 ;
 END
 END vss.gds766
 PIN vss.gds767
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 8.6535 64.214 8.8535 ;
 END
 END vss.gds767
 PIN vss.gds768
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 7.981 63.534 8.181 ;
 END
 END vss.gds768
 PIN vss.gds769
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 8.0595 62.862 8.2595 ;
 END
 END vss.gds769
 PIN vss.gds770
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 8.0595 62.19 8.2595 ;
 END
 END vss.gds770
 PIN vss.gds771
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 8.0595 61.518 8.2595 ;
 END
 END vss.gds771
 PIN vss.gds772
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 8.0595 60.846 8.2595 ;
 END
 END vss.gds772
 PIN vss.gds773
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 7.9635 63.974 8.1635 ;
 END
 END vss.gds773
 PIN vss.gds774
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 8.831 63.746 9.031 ;
 END
 END vss.gds774
 PIN vss.gds775
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 8.0595 64.814 8.2595 ;
 END
 END vss.gds775
 PIN vss.gds776
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 6.458 65.054 6.658 ;
 END
 END vss.gds776
 PIN vss.gds777
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 65.156 10.416 65.212 10.589 ;
 RECT 65.156 6.636 65.212 6.809 ;
 RECT 65.156 7.896 65.212 8.069 ;
 RECT 65.156 9.156 65.212 9.329 ;
 RECT 64.82 9.883 64.876 10.083 ;
 RECT 64.82 8.623 64.876 8.823 ;
 RECT 64.82 7.363 64.876 7.563 ;
 RECT 64.82 6.103 64.876 6.303 ;
 RECT 64.652 7.935 64.708 8.135 ;
 RECT 64.484 7.873 64.54 8.073 ;
 RECT 63.98 7.924 64.036 8.124 ;
 RECT 64.316 7.924 64.372 8.124 ;
 RECT 64.148 7.924 64.204 8.124 ;
 RECT 63.644 7.954 63.7 8.154 ;
 RECT 63.812 7.954 63.868 8.154 ;
 END
 END vss.gds777
 PIN vss.gds778
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 9.018 66.026 9.218 ;
 END
 END vss.gds778
 PIN vss.gds779
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 7.758 66.026 7.958 ;
 END
 END vss.gds779
 PIN vss.gds780
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 6.498 66.026 6.698 ;
 END
 END vss.gds780
 PIN vss.gds781
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 7.213 67.302 7.413 ;
 END
 END vss.gds781
 PIN vss.gds782
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.142 7.843 69.182 8.043 ;
 END
 END vss.gds782
 PIN vss.gds783
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.69 8.0595 69.75 8.2595 ;
 END
 END vss.gds783
 PIN vss.gds784
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.858 8.0595 69.918 8.2595 ;
 END
 END vss.gds784
 PIN vss.gds785
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.194 8.0595 70.254 8.2595 ;
 END
 END vss.gds785
 PIN vss.gds786
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 7.956 66.574 8.156 ;
 END
 END vss.gds786
 PIN vss.gds787
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 8.1 66.318 8.3 ;
 END
 END vss.gds787
 PIN vss.gds788
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 8.0595 70.086 8.2595 ;
 END
 END vss.gds788
 PIN vss.gds789
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 8.0185 68.15 8.2185 ;
 END
 END vss.gds789
 PIN vss.gds790
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 9.733 67.302 9.933 ;
 END
 END vss.gds790
 PIN vss.gds791
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 7.8665 67.646 8.0665 ;
 END
 END vss.gds791
 PIN vss.gds792
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 8.112 67.97 8.312 ;
 END
 END vss.gds792
 PIN vss.gds793
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 5.953 67.302 6.153 ;
 END
 END vss.gds793
 PIN vss.gds794
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 8.473 67.302 8.673 ;
 END
 END vss.gds794
 PIN vss.gds795
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 8.1 65.654 8.3 ;
 END
 END vss.gds795
 PIN vss.gds796
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 8.1 66.998 8.3 ;
 END
 END vss.gds796
 PIN vss.gds797
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 7.9635 68.99 8.1635 ;
 END
 END vss.gds797
 PIN vss.gds798
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.594 8.1155 68.65 8.3155 ;
 END
 END vss.gds798
 PIN vss.gds799
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 7.9635 68.47 8.1635 ;
 END
 END vss.gds799
 PIN vss.gds800
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.522 8.0595 69.582 8.2595 ;
 END
 END vss.gds800
 PIN vss.gds801
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 7.981 69.414 8.181 ;
 END
 END vss.gds801
 PIN vss.gds802
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 67.676 10.436 67.732 10.589 ;
 RECT 65.324 10.389 65.38 10.589 ;
 RECT 66.92 10.433 66.976 10.598 ;
 RECT 66.752 10.433 66.808 10.598 ;
 RECT 65.996 10.433 66.052 10.598 ;
 RECT 65.828 10.433 65.884 10.598 ;
 RECT 66.752 9.4 66.808 9.6 ;
 RECT 67.004 9.403 67.06 9.603 ;
 RECT 67.676 6.656 67.732 6.809 ;
 RECT 65.324 6.609 65.38 6.809 ;
 RECT 66.92 6.653 66.976 6.818 ;
 RECT 66.752 6.653 66.808 6.818 ;
 RECT 65.996 6.653 66.052 6.818 ;
 RECT 65.828 6.653 65.884 6.818 ;
 RECT 67.676 7.916 67.732 8.069 ;
 RECT 65.324 7.869 65.38 8.069 ;
 RECT 66.92 7.913 66.976 8.078 ;
 RECT 66.752 7.913 66.808 8.078 ;
 RECT 65.996 7.913 66.052 8.078 ;
 RECT 65.828 7.913 65.884 8.078 ;
 RECT 67.676 9.176 67.732 9.329 ;
 RECT 65.324 9.129 65.38 9.329 ;
 RECT 66.92 9.173 66.976 9.338 ;
 RECT 66.752 9.173 66.808 9.338 ;
 RECT 65.996 9.173 66.052 9.338 ;
 RECT 65.828 9.173 65.884 9.338 ;
 RECT 65.492 9.749 65.548 9.949 ;
 RECT 65.324 9.749 65.38 9.949 ;
 RECT 66.752 5.62 66.808 5.82 ;
 RECT 67.004 5.623 67.06 5.823 ;
 RECT 66.752 8.14 66.808 8.34 ;
 RECT 67.004 8.143 67.06 8.343 ;
 RECT 66.752 6.88 66.808 7.08 ;
 RECT 67.004 6.883 67.06 7.083 ;
 RECT 68.012 9.8075 68.068 10.0075 ;
 RECT 67.508 10.0595 67.564 10.2595 ;
 RECT 66.164 9.959 66.22 10.159 ;
 RECT 66.584 9.959 66.64 10.159 ;
 RECT 67.508 7.5395 67.564 7.7395 ;
 RECT 68.012 7.2875 68.068 7.4875 ;
 RECT 65.492 7.229 65.548 7.429 ;
 RECT 65.324 7.229 65.38 7.429 ;
 RECT 65.492 5.969 65.548 6.169 ;
 RECT 65.324 5.969 65.38 6.169 ;
 RECT 66.164 6.179 66.22 6.379 ;
 RECT 66.584 6.179 66.64 6.379 ;
 RECT 68.012 8.5475 68.068 8.7475 ;
 RECT 67.508 8.7995 67.564 8.9995 ;
 RECT 66.164 8.699 66.22 8.899 ;
 RECT 66.584 8.699 66.64 8.899 ;
 RECT 65.492 8.489 65.548 8.689 ;
 RECT 65.324 8.489 65.38 8.689 ;
 RECT 66.164 7.439 66.22 7.639 ;
 RECT 66.584 7.439 66.64 7.639 ;
 RECT 67.508 6.2795 67.564 6.4795 ;
 RECT 68.012 6.0275 68.068 6.2275 ;
 RECT 66.332 8.1395 66.388 8.3395 ;
 RECT 69.02 7.954 69.076 8.154 ;
 RECT 68.852 7.9615 68.908 8.1615 ;
 RECT 68.684 7.954 68.74 8.154 ;
 RECT 68.516 7.954 68.572 8.154 ;
 RECT 68.348 7.954 68.404 8.154 ;
 RECT 69.188 7.954 69.244 8.154 ;
 RECT 68.18 8.069 68.236 8.269 ;
 END
 END vss.gds802
 PIN vss.gds803
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.362 8.0595 70.422 8.2595 ;
 END
 END vss.gds803
 PIN vss.gds804
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.53 8.0595 70.59 8.2595 ;
 END
 END vss.gds804
 PIN vss.gds805
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.866 8.0595 70.926 8.2595 ;
 END
 END vss.gds805
 PIN vss.gds806
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.034 8.0595 71.094 8.2595 ;
 END
 END vss.gds806
 PIN vss.gds807
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.202 8.0595 71.262 8.2595 ;
 END
 END vss.gds807
 PIN vss.gds808
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.538 8.0595 71.598 8.2595 ;
 END
 END vss.gds808
 PIN vss.gds809
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.706 8.0595 71.766 8.2595 ;
 END
 END vss.gds809
 PIN vss.gds810
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.874 8.0595 71.934 8.2595 ;
 END
 END vss.gds810
 PIN vss.gds811
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.21 8.0595 72.27 8.2595 ;
 END
 END vss.gds811
 PIN vss.gds812
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.378 8.0595 72.438 8.2595 ;
 END
 END vss.gds812
 PIN vss.gds813
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.546 8.0595 72.606 8.2595 ;
 END
 END vss.gds813
 PIN vss.gds814
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.882 8.0595 72.942 8.2595 ;
 END
 END vss.gds814
 PIN vss.gds815
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.05 8.0595 73.11 8.2595 ;
 END
 END vss.gds815
 PIN vss.gds816
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 8.0595 71.43 8.2595 ;
 END
 END vss.gds816
 PIN vss.gds817
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 8.0595 72.102 8.2595 ;
 END
 END vss.gds817
 PIN vss.gds818
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 8.0595 72.774 8.2595 ;
 END
 END vss.gds818
 PIN vss.gds819
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 8.0595 70.758 8.2595 ;
 END
 END vss.gds819
 PIN vss.gds820
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.554 8.0595 73.614 8.2595 ;
 END
 END vss.gds820
 PIN vss.gds821
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.722 8.0595 73.782 8.2595 ;
 END
 END vss.gds821
 PIN vss.gds822
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.89 8.0595 73.95 8.2595 ;
 END
 END vss.gds822
 PIN vss.gds823
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 8.0595 74.118 8.2595 ;
 END
 END vss.gds823
 PIN vss.gds824
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.394 8.0595 74.454 8.2595 ;
 END
 END vss.gds824
 PIN vss.gds825
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.562 8.0595 74.622 8.2595 ;
 END
 END vss.gds825
 PIN vss.gds826
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 8.0595 74.79 8.2595 ;
 END
 END vss.gds826
 PIN vss.gds827
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.218 8.0595 73.278 8.2595 ;
 END
 END vss.gds827
 PIN vss.gds828
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 8.0595 73.446 8.2595 ;
 END
 END vss.gds828
 PIN vss.gds829
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.226 8.0595 74.286 8.2595 ;
 END
 END vss.gds829
 PIN vss.gds830
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 13.2175 0.29 13.4175 ;
 END
 END vss.gds830
 PIN vss.gds831
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.286 11.741 3.326 11.941 ;
 END
 END vss.gds831
 PIN vss.gds832
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 12.0535 0.602 12.2535 ;
 END
 END vss.gds832
 PIN vss.gds833
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 12.7615 0.942 12.9615 ;
 END
 END vss.gds833
 PIN vss.gds834
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.646 14.2155 1.702 14.4155 ;
 END
 END vss.gds834
 PIN vss.gds835
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 13.4825 1.282 13.6825 ;
 END
 END vss.gds835
 PIN vss.gds836
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 13.7445 2.122 13.9445 ;
 END
 END vss.gds836
 PIN vss.gds837
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.282 12.839 4.338 13.039 ;
 END
 END vss.gds837
 PIN vss.gds838
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 11.346 4.882 11.546 ;
 END
 END vss.gds838
 PIN vss.gds839
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 12.9395 4.194 13.1395 ;
 END
 END vss.gds839
 PIN vss.gds840
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 12.364 5.074 12.564 ;
 END
 END vss.gds840
 PIN vss.gds841
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.746 14.662 2.802 14.862 ;
 END
 END vss.gds841
 PIN vss.gds842
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 15.348 4.882 15.548 ;
 END
 END vss.gds842
 PIN vss.gds843
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 13.4515 4.002 13.6515 ;
 END
 END vss.gds843
 PIN vss.gds844
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 13.5795 5.282 13.7795 ;
 END
 END vss.gds844
 PIN vss.gds845
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.562 15.291 3.602 15.491 ;
 END
 END vss.gds845
 PIN vss.gds846
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 13.8295 2.302 14.0295 ;
 END
 END vss.gds846
 PIN vss.gds847
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 12.8635 3.142 13.0635 ;
 END
 END vss.gds847
 PIN vss.gds848
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 13.356 1.462 13.556 ;
 END
 END vss.gds848
 PIN vss.gds849
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 13.3325 0.718 13.5325 ;
 END
 END vss.gds849
 PIN vss.gds850
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 3.164 14.418 3.22 14.618 ;
 RECT 3.416 14.455 3.472 14.637 ;
 RECT 3.836 14.418 3.892 14.618 ;
 RECT 1.988 14.3475 2.044 14.5475 ;
 RECT 3.5 14.685 3.556 14.836 ;
 RECT 4.004 14.5525 4.06 14.7525 ;
 RECT 3.752 14.685 3.808 14.857 ;
 RECT 0.56 14.7175 0.616 14.9175 ;
 RECT 1.568 14.679 1.624 14.879 ;
 RECT 0.98 14.679 1.036 14.879 ;
 RECT 3.164 13.354 3.22 13.554 ;
 RECT 4.676 13.354 4.732 13.554 ;
 RECT 4.424 13.343 4.48 13.543 ;
 RECT 4.76 10.647 4.816 10.829 ;
 RECT 4.424 10.668 4.48 10.868 ;
 RECT 5.18 10.647 5.236 10.829 ;
 RECT 4.004 10.668 4.06 10.868 ;
 RECT 3.836 10.647 3.892 10.829 ;
 RECT 3.584 10.668 3.64 10.868 ;
 RECT 3.416 10.668 3.472 10.868 ;
 RECT 3.164 12.01 3.22 12.21 ;
 RECT 3.416 11.991 3.472 12.173 ;
 RECT 4.004 12.01 4.06 12.21 ;
 RECT 3.836 12.01 3.892 12.21 ;
 RECT 3.584 11.73 3.64 11.93 ;
 RECT 4.004 11.73 4.06 11.93 ;
 RECT 4.256 11.8645 4.312 12.0645 ;
 RECT 4.76 11.8685 4.816 12.0685 ;
 RECT 4.508 11.8645 4.564 12.0645 ;
 RECT 5.18 11.8685 5.236 12.0685 ;
 RECT 1.568 11.991 1.624 12.191 ;
 RECT 0.98 11.991 1.036 12.191 ;
 RECT 0.56 11.991 0.616 12.191 ;
 RECT 0.56 11.749 0.616 11.949 ;
 RECT 1.568 11.749 1.624 11.949 ;
 RECT 0.98 11.749 1.036 11.949 ;
 RECT 2.156 11.87 2.212 12.07 ;
 RECT 3.164 11.73 3.22 11.93 ;
 RECT 2.66 11.87 2.716 12.07 ;
 RECT 0.56 10.647 0.616 10.847 ;
 RECT 1.568 10.647 1.624 10.847 ;
 RECT 0.98 10.647 1.036 10.847 ;
 RECT 1.904 10.668 1.96 10.868 ;
 RECT 2.156 10.668 2.212 10.868 ;
 RECT 2.408 10.668 2.464 10.868 ;
 RECT 2.912 10.668 2.968 10.868 ;
 RECT 2.66 10.668 2.716 10.868 ;
 RECT 3.164 10.668 3.22 10.868 ;
 RECT 3.164 13.074 3.22 13.274 ;
 RECT 3.416 13.2125 3.472 13.4125 ;
 RECT 4.004 13.214 4.06 13.414 ;
 RECT 3.836 13.214 3.892 13.414 ;
 RECT 4.256 13.2125 4.312 13.4125 ;
 RECT 4.508 13.136 4.564 13.287 ;
 RECT 4.76 13.111 4.816 13.293 ;
 RECT 5.18 13.111 5.236 13.293 ;
 RECT 2.24 13.074 2.296 13.274 ;
 RECT 0.56 13.3735 0.616 13.5735 ;
 RECT 1.568 13.3735 1.624 13.5735 ;
 RECT 0.98 13.3735 1.036 13.5735 ;
 RECT 2.576 13.335 2.632 13.535 ;
 RECT 0.56 13.093 0.616 13.293 ;
 RECT 1.568 13.093 1.624 13.293 ;
 RECT 0.98 13.093 1.036 13.293 ;
 RECT 2.156 13.2605 2.212 13.4605 ;
 RECT 2.912 13.335 2.968 13.535 ;
 RECT 2.744 13.214 2.8 13.414 ;
 RECT 0.56 14.398 0.616 14.598 ;
 RECT 1.568 14.398 1.624 14.598 ;
 RECT 0.98 14.398 1.036 14.598 ;
 RECT 2.492 14.5015 2.548 14.7015 ;
 RECT 2.156 14.558 2.212 14.758 ;
 RECT 2.324 14.5015 2.38 14.7015 ;
 RECT 3.248 14.685 3.304 14.857 ;
 RECT 2.828 14.682 2.884 14.882 ;
 RECT 2.66 14.698 2.716 14.898 ;
 RECT 4.256 14.5565 4.312 14.7565 ;
 RECT 4.676 14.558 4.732 14.758 ;
 RECT 4.424 14.5525 4.48 14.7525 ;
 RECT 1.82 14.398 1.876 14.598 ;
 END
 END vss.gds850
 PIN vss.gds851
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.982 12.105 10.022 12.305 ;
 END
 END vss.gds851
 PIN vss.gds852
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.31 12.105 9.35 12.305 ;
 END
 END vss.gds852
 PIN vss.gds853
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.638 12.105 8.678 12.305 ;
 END
 END vss.gds853
 PIN vss.gds854
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.966 12.105 8.006 12.305 ;
 END
 END vss.gds854
 PIN vss.gds855
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.294 12.105 7.334 12.305 ;
 END
 END vss.gds855
 PIN vss.gds856
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.778 12.41 9.824 12.61 ;
 END
 END vss.gds856
 PIN vss.gds857
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.174 12.5875 10.214 12.7875 ;
 END
 END vss.gds857
 PIN vss.gds858
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.106 12.41 9.152 12.61 ;
 END
 END vss.gds858
 PIN vss.gds859
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.502 12.5875 9.542 12.7875 ;
 END
 END vss.gds859
 PIN vss.gds860
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.434 12.41 8.48 12.61 ;
 END
 END vss.gds860
 PIN vss.gds861
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.762 12.41 7.808 12.61 ;
 END
 END vss.gds861
 PIN vss.gds862
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.09 12.41 7.136 12.61 ;
 END
 END vss.gds862
 PIN vss.gds863
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.83 12.5875 8.87 12.7875 ;
 END
 END vss.gds863
 PIN vss.gds864
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.158 12.5875 8.198 12.7875 ;
 END
 END vss.gds864
 PIN vss.gds865
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.486 12.5875 7.526 12.7875 ;
 END
 END vss.gds865
 PIN vss.gds866
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 13.1145 9.69 13.3145 ;
 END
 END vss.gds866
 PIN vss.gds867
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 13.1145 8.346 13.3145 ;
 END
 END vss.gds867
 PIN vss.gds868
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 13.1145 9.018 13.3145 ;
 END
 END vss.gds868
 PIN vss.gds869
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.942 13.1145 7.002 13.3145 ;
 END
 END vss.gds869
 PIN vss.gds870
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 13.1145 7.674 13.3145 ;
 END
 END vss.gds870
 PIN vss.gds871
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 13.45 5.474 13.65 ;
 END
 END vss.gds871
 PIN vss.gds872
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 13.9715 5.986 14.1715 ;
 END
 END vss.gds872
 PIN vss.gds873
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.734 13.7955 6.774 13.9955 ;
 END
 END vss.gds873
 PIN vss.gds874
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.606 13.6715 6.646 13.8715 ;
 END
 END vss.gds874
 PIN vss.gds875
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 13.838 5.73 14.038 ;
 END
 END vss.gds875
 PIN vss.gds876
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 13.031 6.434 13.231 ;
 END
 END vss.gds876
 PIN vss.gds877
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 11.31 6.178 11.51 ;
 END
 END vss.gds877
 PIN vss.gds878
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 5.432 13.354 5.488 13.554 ;
 RECT 5.6 13.354 5.656 13.554 ;
 RECT 5.768 13.354 5.824 13.554 ;
 RECT 5.936 13.354 5.992 13.554 ;
 RECT 6.104 13.354 6.16 13.554 ;
 RECT 6.272 10.668 6.328 10.868 ;
 RECT 6.104 10.668 6.16 10.868 ;
 RECT 5.852 10.668 5.908 10.868 ;
 RECT 5.684 10.668 5.74 10.868 ;
 RECT 9.968 11.11 10.024 11.31 ;
 RECT 9.8 11.11 9.856 11.31 ;
 RECT 10.136 11.11 10.192 11.31 ;
 RECT 9.296 11.11 9.352 11.31 ;
 RECT 9.128 11.11 9.184 11.31 ;
 RECT 9.464 11.11 9.52 11.31 ;
 RECT 9.632 11.101 9.688 11.301 ;
 RECT 8.624 11.11 8.68 11.31 ;
 RECT 8.456 11.11 8.512 11.31 ;
 RECT 8.792 11.11 8.848 11.31 ;
 RECT 8.96 11.101 9.016 11.301 ;
 RECT 7.952 11.11 8.008 11.31 ;
 RECT 7.784 11.11 7.84 11.31 ;
 RECT 8.12 11.11 8.176 11.31 ;
 RECT 8.288 11.101 8.344 11.301 ;
 RECT 6.944 11.101 7 11.301 ;
 RECT 7.28 11.11 7.336 11.31 ;
 RECT 7.112 11.11 7.168 11.31 ;
 RECT 7.448 11.11 7.504 11.31 ;
 RECT 7.616 11.101 7.672 11.301 ;
 RECT 9.632 14.4275 9.688 14.6275 ;
 RECT 8.96 14.4275 9.016 14.6275 ;
 RECT 8.288 14.4275 8.344 14.6275 ;
 RECT 6.944 14.222 7 14.422 ;
 RECT 7.616 14.4275 7.672 14.6275 ;
 RECT 6.272 11.87 6.328 12.07 ;
 RECT 6.104 11.87 6.16 12.07 ;
 RECT 5.852 11.87 5.908 12.07 ;
 RECT 5.684 11.87 5.74 12.07 ;
 RECT 6.44 11.73 6.496 11.93 ;
 RECT 6.44 12.01 6.496 12.21 ;
 RECT 9.968 12.6525 10.024 12.8525 ;
 RECT 9.8 12.6525 9.856 12.8525 ;
 RECT 10.136 12.6525 10.192 12.8525 ;
 RECT 9.296 12.6525 9.352 12.8525 ;
 RECT 9.128 12.6525 9.184 12.8525 ;
 RECT 9.632 12.6525 9.688 12.8525 ;
 RECT 9.464 12.6525 9.52 12.8525 ;
 RECT 8.624 12.6525 8.68 12.8525 ;
 RECT 8.456 12.6525 8.512 12.8525 ;
 RECT 8.96 12.6525 9.016 12.8525 ;
 RECT 8.792 12.6525 8.848 12.8525 ;
 RECT 7.952 12.6525 8.008 12.8525 ;
 RECT 7.784 12.6525 7.84 12.8525 ;
 RECT 8.288 12.6525 8.344 12.8525 ;
 RECT 8.12 12.6525 8.176 12.8525 ;
 RECT 7.28 12.6525 7.336 12.8525 ;
 RECT 6.944 12.6525 7 12.8525 ;
 RECT 7.112 12.6525 7.168 12.8525 ;
 RECT 7.616 12.6525 7.672 12.8525 ;
 RECT 7.448 12.6525 7.504 12.8525 ;
 RECT 6.44 10.668 6.496 10.868 ;
 RECT 6.104 13.074 6.16 13.274 ;
 RECT 5.852 13.074 5.908 13.274 ;
 RECT 5.684 13.074 5.74 13.274 ;
 RECT 6.44 13.214 6.496 13.414 ;
 RECT 6.272 13.214 6.328 13.414 ;
 RECT 5.432 14.558 5.488 14.758 ;
 RECT 5.6 14.558 5.656 14.758 ;
 RECT 5.768 14.558 5.824 14.758 ;
 RECT 5.936 14.558 5.992 14.758 ;
 RECT 6.44 14.558 6.496 14.758 ;
 RECT 6.104 14.558 6.16 14.758 ;
 RECT 6.272 14.558 6.328 14.758 ;
 END
 END vss.gds878
 PIN vss.gds879
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.998 12.105 12.038 12.305 ;
 END
 END vss.gds879
 PIN vss.gds880
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.326 12.105 11.366 12.305 ;
 END
 END vss.gds880
 PIN vss.gds881
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.654 12.105 10.694 12.305 ;
 END
 END vss.gds881
 PIN vss.gds882
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.794 12.41 11.84 12.61 ;
 END
 END vss.gds882
 PIN vss.gds883
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.19 12.5875 12.23 12.7875 ;
 END
 END vss.gds883
 PIN vss.gds884
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.122 12.41 11.168 12.61 ;
 END
 END vss.gds884
 PIN vss.gds885
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.518 12.5875 11.558 12.7875 ;
 END
 END vss.gds885
 PIN vss.gds886
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.45 12.41 10.496 12.61 ;
 END
 END vss.gds886
 PIN vss.gds887
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.846 12.5875 10.886 12.7875 ;
 END
 END vss.gds887
 PIN vss.gds888
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.262 11.488 14.318 11.688 ;
 END
 END vss.gds888
 PIN vss.gds889
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 11.699 14.87 11.899 ;
 END
 END vss.gds889
 PIN vss.gds890
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.422 11.5435 13.478 11.7435 ;
 END
 END vss.gds890
 PIN vss.gds891
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 12.961 13.658 13.161 ;
 END
 END vss.gds891
 PIN vss.gds892
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 13.1145 11.706 13.3145 ;
 END
 END vss.gds892
 PIN vss.gds893
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 13.1145 11.034 13.3145 ;
 END
 END vss.gds893
 PIN vss.gds894
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 13.0485 15.162 13.2485 ;
 END
 END vss.gds894
 PIN vss.gds895
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 13.1145 10.362 13.3145 ;
 END
 END vss.gds895
 PIN vss.gds896
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 13.031 14.498 13.231 ;
 END
 END vss.gds896
 PIN vss.gds897
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 12.961 12.818 13.161 ;
 END
 END vss.gds897
 PIN vss.gds898
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 12.9745 12.378 13.1745 ;
 END
 END vss.gds898
 PIN vss.gds899
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 13.406 12.59 13.606 ;
 END
 END vss.gds899
 PIN vss.gds900
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 11.8645 13.058 12.0645 ;
 END
 END vss.gds900
 PIN vss.gds901
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 12.74 14.698 12.796 14.898 ;
 RECT 14.252 14.679 14.308 14.861 ;
 RECT 15.092 14.739 15.148 14.939 ;
 RECT 14.756 14.698 14.812 14.898 ;
 RECT 14.504 14.679 14.56 14.861 ;
 RECT 13.496 13.354 13.552 13.554 ;
 RECT 14.336 13.354 14.392 13.554 ;
 RECT 13.916 13.354 13.972 13.554 ;
 RECT 14.672 13.335 14.728 13.517 ;
 RECT 14.84 13.354 14.896 13.554 ;
 RECT 13.58 10.668 13.636 10.868 ;
 RECT 12.908 10.668 12.964 10.868 ;
 RECT 13.916 10.668 13.972 10.868 ;
 RECT 14.252 10.668 14.308 10.868 ;
 RECT 14.588 10.668 14.644 10.868 ;
 RECT 14.924 10.668 14.98 10.868 ;
 RECT 12.656 12.01 12.712 12.21 ;
 RECT 13.244 11.991 13.3 12.173 ;
 RECT 12.656 11.73 12.712 11.93 ;
 RECT 13.244 11.767 13.3 11.949 ;
 RECT 13.916 11.87 13.972 12.07 ;
 RECT 13.076 13.4245 13.132 13.6245 ;
 RECT 13.328 13.4245 13.384 13.6245 ;
 RECT 14.168 13.4245 14.224 13.6245 ;
 RECT 13.748 13.4245 13.804 13.6245 ;
 RECT 15.176 13.4245 15.232 13.6245 ;
 RECT 13.244 14.558 13.3 14.758 ;
 RECT 14.252 14.455 14.308 14.637 ;
 RECT 13.916 14.558 13.972 14.758 ;
 RECT 15.092 14.418 15.148 14.618 ;
 RECT 14.756 14.418 14.812 14.618 ;
 RECT 14.588 14.455 14.644 14.637 ;
 RECT 13.244 10.629 13.3 10.829 ;
 RECT 11.984 11.11 12.04 11.31 ;
 RECT 11.816 11.11 11.872 11.31 ;
 RECT 12.152 11.11 12.208 11.31 ;
 RECT 12.32 11.101 12.376 11.301 ;
 RECT 11.312 11.11 11.368 11.31 ;
 RECT 11.144 11.11 11.2 11.31 ;
 RECT 11.48 11.11 11.536 11.31 ;
 RECT 11.648 11.101 11.704 11.301 ;
 RECT 10.64 11.11 10.696 11.31 ;
 RECT 10.472 11.11 10.528 11.31 ;
 RECT 10.808 11.11 10.864 11.31 ;
 RECT 10.976 11.101 11.032 11.301 ;
 RECT 10.304 11.101 10.36 11.301 ;
 RECT 12.32 14.4275 12.376 14.6275 ;
 RECT 11.648 14.4275 11.704 14.6275 ;
 RECT 10.976 14.4275 11.032 14.6275 ;
 RECT 10.304 14.4275 10.36 14.6275 ;
 RECT 12.824 10.474 12.88 10.674 ;
 RECT 11.984 12.6525 12.04 12.8525 ;
 RECT 11.816 12.6525 11.872 12.8525 ;
 RECT 12.32 12.6525 12.376 12.8525 ;
 RECT 12.152 12.6525 12.208 12.8525 ;
 RECT 11.312 12.6525 11.368 12.8525 ;
 RECT 11.144 12.6525 11.2 12.8525 ;
 RECT 11.648 12.6525 11.704 12.8525 ;
 RECT 11.48 12.6525 11.536 12.8525 ;
 RECT 10.64 12.6525 10.696 12.8525 ;
 RECT 10.472 12.6525 10.528 12.8525 ;
 RECT 10.976 12.6525 11.032 12.8525 ;
 RECT 10.808 12.6525 10.864 12.8525 ;
 RECT 10.304 12.6525 10.36 12.8525 ;
 RECT 13.328 10.474 13.384 10.674 ;
 RECT 13.16 10.474 13.216 10.674 ;
 RECT 12.488 10.474 12.544 10.674 ;
 RECT 12.992 10.474 13.048 10.674 ;
 RECT 12.656 10.5945 12.712 10.7945 ;
 RECT 13.496 13.074 13.552 13.274 ;
 RECT 13.076 13.074 13.132 13.274 ;
 RECT 13.916 13.074 13.972 13.274 ;
 RECT 14.336 13.074 14.392 13.274 ;
 RECT 14.84 13.074 14.896 13.274 ;
 RECT 14.672 13.111 14.728 13.293 ;
 RECT 15.176 13.0035 15.232 13.2035 ;
 END
 END vss.gds901
 PIN vss.gds902
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.894 12.105 19.934 12.305 ;
 END
 END vss.gds902
 PIN vss.gds903
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.222 12.105 19.262 12.305 ;
 END
 END vss.gds903
 PIN vss.gds904
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.69 12.41 19.736 12.61 ;
 END
 END vss.gds904
 PIN vss.gds905
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.086 12.5875 20.126 12.7875 ;
 END
 END vss.gds905
 PIN vss.gds906
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.018 12.41 19.064 12.61 ;
 END
 END vss.gds906
 PIN vss.gds907
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.414 12.5875 19.454 12.7875 ;
 END
 END vss.gds907
 PIN vss.gds908
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.346 12.41 18.392 12.61 ;
 END
 END vss.gds908
 PIN vss.gds909
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.742 12.5875 18.782 12.7875 ;
 END
 END vss.gds909
 PIN vss.gds910
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.594 14.951 16.65 15.151 ;
 END
 END vss.gds910
 PIN vss.gds911
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 13.1145 20.274 13.3145 ;
 END
 END vss.gds911
 PIN vss.gds912
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 13.1445 16.146 13.3445 ;
 END
 END vss.gds912
 PIN vss.gds913
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.598 13.515 17.654 13.715 ;
 END
 END vss.gds913
 PIN vss.gds914
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.17 14.5535 16.226 14.7535 ;
 END
 END vss.gds914
 PIN vss.gds915
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 14.29 17.314 14.49 ;
 END
 END vss.gds915
 PIN vss.gds916
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 11.346 16.814 11.546 ;
 END
 END vss.gds916
 PIN vss.gds917
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 11.488 15.418 11.688 ;
 END
 END vss.gds917
 PIN vss.gds918
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.55 12.105 18.59 12.305 ;
 END
 END vss.gds918
 PIN vss.gds919
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 13.1145 19.602 13.3145 ;
 END
 END vss.gds919
 PIN vss.gds920
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 13.1145 18.93 13.3145 ;
 END
 END vss.gds920
 PIN vss.gds921
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 13.1495 16.994 13.3495 ;
 END
 END vss.gds921
 PIN vss.gds922
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 13.347 15.842 13.547 ;
 END
 END vss.gds922
 PIN vss.gds923
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 13.1955 17.834 13.3955 ;
 END
 END vss.gds923
 PIN vss.gds924
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 13.048 16.49 13.248 ;
 END
 END vss.gds924
 PIN vss.gds925
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 13.1145 18.258 13.3145 ;
 END
 END vss.gds925
 PIN vss.gds926
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 10.877 17.314 11.077 ;
 END
 END vss.gds926
 PIN vss.gds927
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 15.428 14.698 15.484 14.898 ;
 RECT 16.016 14.698 16.072 14.898 ;
 RECT 15.848 14.698 15.904 14.898 ;
 RECT 16.52 14.679 16.576 14.861 ;
 RECT 16.268 14.679 16.324 14.861 ;
 RECT 17.108 14.698 17.164 14.898 ;
 RECT 17.276 14.698 17.332 14.898 ;
 RECT 16.1 13.335 16.156 13.513 ;
 RECT 15.512 13.354 15.568 13.554 ;
 RECT 15.848 13.335 15.904 13.513 ;
 RECT 16.604 13.354 16.66 13.554 ;
 RECT 17.108 13.354 17.164 13.554 ;
 RECT 17.528 13.354 17.584 13.554 ;
 RECT 15.932 10.668 15.988 10.868 ;
 RECT 16.268 10.668 16.324 10.868 ;
 RECT 16.604 10.668 16.66 10.868 ;
 RECT 16.94 10.668 16.996 10.868 ;
 RECT 15.932 12.01 15.988 12.21 ;
 RECT 15.764 12.01 15.82 12.21 ;
 RECT 15.596 12.01 15.652 12.21 ;
 RECT 15.428 12.01 15.484 12.21 ;
 RECT 16.604 12.01 16.66 12.21 ;
 RECT 16.184 11.992 16.24 12.169 ;
 RECT 15.932 11.73 15.988 11.93 ;
 RECT 15.764 11.73 15.82 11.93 ;
 RECT 15.596 11.73 15.652 11.93 ;
 RECT 15.428 11.73 15.484 11.93 ;
 RECT 16.184 11.771 16.24 11.949 ;
 RECT 16.352 11.767 16.408 11.967 ;
 RECT 16.688 11.73 16.744 11.93 ;
 RECT 18.2 14.222 18.256 14.422 ;
 RECT 19.88 11.11 19.936 11.31 ;
 RECT 19.712 11.11 19.768 11.31 ;
 RECT 20.048 11.11 20.104 11.31 ;
 RECT 20.216 11.101 20.272 11.301 ;
 RECT 19.208 11.11 19.264 11.31 ;
 RECT 19.04 11.11 19.096 11.31 ;
 RECT 19.376 11.11 19.432 11.31 ;
 RECT 19.544 11.101 19.6 11.301 ;
 RECT 18.2 11.101 18.256 11.301 ;
 RECT 17.276 10.629 17.332 10.829 ;
 RECT 18.536 11.11 18.592 11.31 ;
 RECT 18.368 11.11 18.424 11.31 ;
 RECT 18.704 11.11 18.76 11.31 ;
 RECT 18.872 11.101 18.928 11.301 ;
 RECT 17.78 14.7685 17.836 14.9685 ;
 RECT 16.1 14.455 16.156 14.637 ;
 RECT 15.428 14.418 15.484 14.618 ;
 RECT 15.764 14.455 15.82 14.637 ;
 RECT 16.604 14.418 16.66 14.618 ;
 RECT 17.192 14.455 17.248 14.637 ;
 RECT 20.216 14.4275 20.272 14.6275 ;
 RECT 19.544 14.4275 19.6 14.6275 ;
 RECT 18.872 14.4275 18.928 14.6275 ;
 RECT 17.864 10.526 17.92 10.726 ;
 RECT 17.696 10.474 17.752 10.674 ;
 RECT 17.528 10.474 17.584 10.674 ;
 RECT 17.36 10.526 17.416 10.726 ;
 RECT 17.192 10.474 17.248 10.674 ;
 RECT 17.528 11.9815 17.584 12.1815 ;
 RECT 16.94 11.87 16.996 12.07 ;
 RECT 17.276 11.87 17.332 12.07 ;
 RECT 17.108 11.87 17.164 12.07 ;
 RECT 17.864 11.73 17.92 11.93 ;
 RECT 17.78 12.051 17.836 12.251 ;
 RECT 19.88 12.6525 19.936 12.8525 ;
 RECT 19.712 12.6525 19.768 12.8525 ;
 RECT 20.216 12.6525 20.272 12.8525 ;
 RECT 20.048 12.6525 20.104 12.8525 ;
 RECT 19.208 12.6525 19.264 12.8525 ;
 RECT 19.04 12.6525 19.096 12.8525 ;
 RECT 19.544 12.6525 19.6 12.8525 ;
 RECT 19.376 12.6525 19.432 12.8525 ;
 RECT 18.536 12.6525 18.592 12.8525 ;
 RECT 18.2 12.6525 18.256 12.8525 ;
 RECT 18.368 12.6525 18.424 12.8525 ;
 RECT 18.872 12.6525 18.928 12.8525 ;
 RECT 18.704 12.6525 18.76 12.8525 ;
 RECT 18.032 10.474 18.088 10.674 ;
 RECT 16.1 13.115 16.156 13.287 ;
 RECT 15.848 13.115 15.904 13.287 ;
 RECT 15.512 13.074 15.568 13.274 ;
 RECT 16.52 13.074 16.576 13.274 ;
 RECT 17.528 13.074 17.584 13.274 ;
 RECT 17.024 13.074 17.08 13.274 ;
 END
 END vss.gds927
 PIN vss.gds928
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.018 12.105 25.058 12.305 ;
 END
 END vss.gds928
 PIN vss.gds929
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.346 12.105 24.386 12.305 ;
 END
 END vss.gds929
 PIN vss.gds930
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.254 12.105 23.294 12.305 ;
 END
 END vss.gds930
 PIN vss.gds931
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.582 12.105 22.622 12.305 ;
 END
 END vss.gds931
 PIN vss.gds932
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.91 12.105 21.95 12.305 ;
 END
 END vss.gds932
 PIN vss.gds933
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.238 12.105 21.278 12.305 ;
 END
 END vss.gds933
 PIN vss.gds934
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.566 12.105 20.606 12.305 ;
 END
 END vss.gds934
 PIN vss.gds935
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.814 12.41 24.86 12.61 ;
 END
 END vss.gds935
 PIN vss.gds936
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.21 12.5875 25.25 12.7875 ;
 END
 END vss.gds936
 PIN vss.gds937
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.142 12.41 24.188 12.61 ;
 END
 END vss.gds937
 PIN vss.gds938
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.538 12.5875 24.578 12.7875 ;
 END
 END vss.gds938
 PIN vss.gds939
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.05 12.41 23.096 12.61 ;
 END
 END vss.gds939
 PIN vss.gds940
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.446 12.5875 23.486 12.7875 ;
 END
 END vss.gds940
 PIN vss.gds941
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.378 12.41 22.424 12.61 ;
 END
 END vss.gds941
 PIN vss.gds942
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.774 12.5875 22.814 12.7875 ;
 END
 END vss.gds942
 PIN vss.gds943
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.706 12.41 21.752 12.61 ;
 END
 END vss.gds943
 PIN vss.gds944
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.102 12.5875 22.142 12.7875 ;
 END
 END vss.gds944
 PIN vss.gds945
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.034 12.41 21.08 12.61 ;
 END
 END vss.gds945
 PIN vss.gds946
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.43 12.5875 21.47 12.7875 ;
 END
 END vss.gds946
 PIN vss.gds947
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.362 12.41 20.408 12.61 ;
 END
 END vss.gds947
 PIN vss.gds948
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.758 12.5875 20.798 12.7875 ;
 END
 END vss.gds948
 PIN vss.gds949
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 13.1145 24.726 13.3145 ;
 END
 END vss.gds949
 PIN vss.gds950
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 13.1145 22.962 13.3145 ;
 END
 END vss.gds950
 PIN vss.gds951
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 13.1145 22.29 13.3145 ;
 END
 END vss.gds951
 PIN vss.gds952
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 13.1145 21.618 13.3145 ;
 END
 END vss.gds952
 PIN vss.gds953
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 13.1145 20.946 13.3145 ;
 END
 END vss.gds953
 PIN vss.gds954
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.994 13.1765 24.054 13.3765 ;
 END
 END vss.gds954
 PIN vss.gds955
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.722 13.852 23.762 14.052 ;
 END
 END vss.gds955
 PIN vss.gds956
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.866 13.852 23.906 14.052 ;
 END
 END vss.gds956
 PIN vss.gds957
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 13.1765 23.634 13.3765 ;
 END
 END vss.gds957
 PIN vss.gds958
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 23.996 14.222 24.052 14.422 ;
 RECT 25.004 11.11 25.06 11.31 ;
 RECT 24.836 11.11 24.892 11.31 ;
 RECT 25.172 11.11 25.228 11.31 ;
 RECT 24.668 11.101 24.724 11.301 ;
 RECT 23.996 10.9305 24.052 11.1305 ;
 RECT 24.332 11.11 24.388 11.31 ;
 RECT 24.164 11.11 24.22 11.31 ;
 RECT 24.5 11.11 24.556 11.31 ;
 RECT 23.24 11.11 23.296 11.31 ;
 RECT 23.072 11.11 23.128 11.31 ;
 RECT 23.408 11.11 23.464 11.31 ;
 RECT 23.576 11.101 23.632 11.301 ;
 RECT 22.568 11.11 22.624 11.31 ;
 RECT 22.4 11.11 22.456 11.31 ;
 RECT 22.736 11.11 22.792 11.31 ;
 RECT 22.904 11.101 22.96 11.301 ;
 RECT 21.896 11.11 21.952 11.31 ;
 RECT 21.728 11.11 21.784 11.31 ;
 RECT 22.064 11.11 22.12 11.31 ;
 RECT 22.232 11.101 22.288 11.301 ;
 RECT 21.224 11.11 21.28 11.31 ;
 RECT 21.056 11.11 21.112 11.31 ;
 RECT 21.392 11.11 21.448 11.31 ;
 RECT 21.56 11.101 21.616 11.301 ;
 RECT 20.888 11.101 20.944 11.301 ;
 RECT 20.552 11.11 20.608 11.31 ;
 RECT 20.72 11.11 20.776 11.31 ;
 RECT 20.384 11.11 20.44 11.31 ;
 RECT 24.668 14.4275 24.724 14.6275 ;
 RECT 23.576 14.4275 23.632 14.6275 ;
 RECT 22.904 14.4275 22.96 14.6275 ;
 RECT 22.232 14.4275 22.288 14.6275 ;
 RECT 21.56 14.4275 21.616 14.6275 ;
 RECT 20.888 14.4275 20.944 14.6275 ;
 RECT 25.004 12.6525 25.06 12.8525 ;
 RECT 24.836 12.6525 24.892 12.8525 ;
 RECT 25.172 12.6525 25.228 12.8525 ;
 RECT 24.332 12.6525 24.388 12.8525 ;
 RECT 23.996 12.6525 24.052 12.8525 ;
 RECT 24.164 12.6525 24.22 12.8525 ;
 RECT 24.668 12.6525 24.724 12.8525 ;
 RECT 24.5 12.6525 24.556 12.8525 ;
 RECT 23.24 12.6525 23.296 12.8525 ;
 RECT 23.072 12.6525 23.128 12.8525 ;
 RECT 23.576 12.6525 23.632 12.8525 ;
 RECT 23.408 12.6525 23.464 12.8525 ;
 RECT 22.568 12.6525 22.624 12.8525 ;
 RECT 22.4 12.6525 22.456 12.8525 ;
 RECT 22.904 12.6525 22.96 12.8525 ;
 RECT 22.736 12.6525 22.792 12.8525 ;
 RECT 21.896 12.6525 21.952 12.8525 ;
 RECT 21.728 12.6525 21.784 12.8525 ;
 RECT 22.232 12.6525 22.288 12.8525 ;
 RECT 22.064 12.6525 22.12 12.8525 ;
 RECT 21.224 12.6525 21.28 12.8525 ;
 RECT 21.056 12.6525 21.112 12.8525 ;
 RECT 21.56 12.6525 21.616 12.8525 ;
 RECT 21.392 12.6525 21.448 12.8525 ;
 RECT 20.552 12.6525 20.608 12.8525 ;
 RECT 20.888 12.6525 20.944 12.8525 ;
 RECT 20.72 12.6525 20.776 12.8525 ;
 RECT 20.384 12.6525 20.44 12.8525 ;
 RECT 23.744 12.812 23.8 13.012 ;
 END
 END vss.gds958
 PIN vss.gds959
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.05 12.105 29.09 12.305 ;
 END
 END vss.gds959
 PIN vss.gds960
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.378 12.105 28.418 12.305 ;
 END
 END vss.gds960
 PIN vss.gds961
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.706 12.105 27.746 12.305 ;
 END
 END vss.gds961
 PIN vss.gds962
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.034 12.105 27.074 12.305 ;
 END
 END vss.gds962
 PIN vss.gds963
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.362 12.105 26.402 12.305 ;
 END
 END vss.gds963
 PIN vss.gds964
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.69 12.105 25.73 12.305 ;
 END
 END vss.gds964
 PIN vss.gds965
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.846 12.41 28.892 12.61 ;
 END
 END vss.gds965
 PIN vss.gds966
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.242 12.5875 29.282 12.7875 ;
 END
 END vss.gds966
 PIN vss.gds967
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.174 12.41 28.22 12.61 ;
 END
 END vss.gds967
 PIN vss.gds968
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.57 12.5875 28.61 12.7875 ;
 END
 END vss.gds968
 PIN vss.gds969
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.502 12.41 27.548 12.61 ;
 END
 END vss.gds969
 PIN vss.gds970
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.898 12.5875 27.938 12.7875 ;
 END
 END vss.gds970
 PIN vss.gds971
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.83 12.41 26.876 12.61 ;
 END
 END vss.gds971
 PIN vss.gds972
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.226 12.5875 27.266 12.7875 ;
 END
 END vss.gds972
 PIN vss.gds973
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.158 12.41 26.204 12.61 ;
 END
 END vss.gds973
 PIN vss.gds974
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.554 12.5875 26.594 12.7875 ;
 END
 END vss.gds974
 PIN vss.gds975
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.486 12.41 25.532 12.61 ;
 END
 END vss.gds975
 PIN vss.gds976
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.882 12.5875 25.922 12.7875 ;
 END
 END vss.gds976
 PIN vss.gds977
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 11.8645 30.11 12.0645 ;
 END
 END vss.gds977
 PIN vss.gds978
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 12.9745 29.43 13.1745 ;
 END
 END vss.gds978
 PIN vss.gds979
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 13.1145 28.758 13.3145 ;
 END
 END vss.gds979
 PIN vss.gds980
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 13.1145 28.086 13.3145 ;
 END
 END vss.gds980
 PIN vss.gds981
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 13.1145 27.414 13.3145 ;
 END
 END vss.gds981
 PIN vss.gds982
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 13.1145 26.742 13.3145 ;
 END
 END vss.gds982
 PIN vss.gds983
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 13.1145 26.07 13.3145 ;
 END
 END vss.gds983
 PIN vss.gds984
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 13.1145 25.398 13.3145 ;
 END
 END vss.gds984
 PIN vss.gds985
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 12.961 29.87 13.161 ;
 END
 END vss.gds985
 PIN vss.gds986
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 13.406 29.642 13.606 ;
 END
 END vss.gds986
 PIN vss.gds987
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.792 14.698 29.848 14.898 ;
 RECT 30.128 13.074 30.184 13.274 ;
 RECT 29.96 10.668 30.016 10.868 ;
 RECT 29.708 12.01 29.764 12.21 ;
 RECT 29.708 11.73 29.764 11.93 ;
 RECT 30.128 13.4245 30.184 13.6245 ;
 RECT 29.036 11.11 29.092 11.31 ;
 RECT 28.868 11.11 28.924 11.31 ;
 RECT 29.204 11.11 29.26 11.31 ;
 RECT 29.372 11.101 29.428 11.301 ;
 RECT 28.364 11.11 28.42 11.31 ;
 RECT 28.196 11.11 28.252 11.31 ;
 RECT 28.532 11.11 28.588 11.31 ;
 RECT 28.7 11.101 28.756 11.301 ;
 RECT 27.692 11.11 27.748 11.31 ;
 RECT 27.524 11.11 27.58 11.31 ;
 RECT 27.86 11.11 27.916 11.31 ;
 RECT 28.028 11.101 28.084 11.301 ;
 RECT 27.02 11.11 27.076 11.31 ;
 RECT 26.852 11.11 26.908 11.31 ;
 RECT 27.188 11.11 27.244 11.31 ;
 RECT 27.356 11.101 27.412 11.301 ;
 RECT 26.348 11.11 26.404 11.31 ;
 RECT 26.18 11.11 26.236 11.31 ;
 RECT 26.516 11.11 26.572 11.31 ;
 RECT 26.684 11.101 26.74 11.301 ;
 RECT 25.676 11.11 25.732 11.31 ;
 RECT 25.508 11.11 25.564 11.31 ;
 RECT 25.844 11.11 25.9 11.31 ;
 RECT 26.012 11.101 26.068 11.301 ;
 RECT 25.34 11.101 25.396 11.301 ;
 RECT 29.372 14.4275 29.428 14.6275 ;
 RECT 28.7 14.4275 28.756 14.6275 ;
 RECT 28.028 14.4275 28.084 14.6275 ;
 RECT 27.356 14.4275 27.412 14.6275 ;
 RECT 26.684 14.4275 26.74 14.6275 ;
 RECT 26.012 14.4275 26.068 14.6275 ;
 RECT 25.34 14.4275 25.396 14.6275 ;
 RECT 29.876 10.474 29.932 10.674 ;
 RECT 29.54 10.474 29.596 10.674 ;
 RECT 30.212 10.474 30.268 10.674 ;
 RECT 30.044 10.474 30.1 10.674 ;
 RECT 29.708 10.5945 29.764 10.7945 ;
 RECT 29.036 12.6525 29.092 12.8525 ;
 RECT 28.868 12.6525 28.924 12.8525 ;
 RECT 29.372 12.6525 29.428 12.8525 ;
 RECT 29.204 12.6525 29.26 12.8525 ;
 RECT 28.364 12.6525 28.42 12.8525 ;
 RECT 28.196 12.6525 28.252 12.8525 ;
 RECT 28.7 12.6525 28.756 12.8525 ;
 RECT 28.532 12.6525 28.588 12.8525 ;
 RECT 27.692 12.6525 27.748 12.8525 ;
 RECT 27.524 12.6525 27.58 12.8525 ;
 RECT 28.028 12.6525 28.084 12.8525 ;
 RECT 27.86 12.6525 27.916 12.8525 ;
 RECT 27.02 12.6525 27.076 12.8525 ;
 RECT 26.852 12.6525 26.908 12.8525 ;
 RECT 27.356 12.6525 27.412 12.8525 ;
 RECT 27.188 12.6525 27.244 12.8525 ;
 RECT 26.348 12.6525 26.404 12.8525 ;
 RECT 26.18 12.6525 26.236 12.8525 ;
 RECT 26.684 12.6525 26.74 12.8525 ;
 RECT 26.516 12.6525 26.572 12.8525 ;
 RECT 25.676 12.6525 25.732 12.8525 ;
 RECT 25.508 12.6525 25.564 12.8525 ;
 RECT 26.012 12.6525 26.068 12.8525 ;
 RECT 25.844 12.6525 25.9 12.8525 ;
 RECT 25.34 12.6525 25.396 12.8525 ;
 END
 END vss.gds987
 PIN vss.gds988
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.646 14.951 33.702 15.151 ;
 END
 END vss.gds988
 PIN vss.gds989
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.222 14.5535 33.278 14.7535 ;
 END
 END vss.gds989
 PIN vss.gds990
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 13.1445 33.198 13.3445 ;
 END
 END vss.gds990
 PIN vss.gds991
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 14.29 34.366 14.49 ;
 END
 END vss.gds991
 PIN vss.gds992
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.474 11.5435 30.53 11.7435 ;
 END
 END vss.gds992
 PIN vss.gds993
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 13.347 32.894 13.547 ;
 END
 END vss.gds993
 PIN vss.gds994
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.65 13.515 34.706 13.715 ;
 END
 END vss.gds994
 PIN vss.gds995
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.314 11.488 31.37 11.688 ;
 END
 END vss.gds995
 PIN vss.gds996
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 13.0485 32.214 13.2485 ;
 END
 END vss.gds996
 PIN vss.gds997
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 11.699 31.922 11.899 ;
 END
 END vss.gds997
 PIN vss.gds998
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 11.488 32.47 11.688 ;
 END
 END vss.gds998
 PIN vss.gds999
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 12.961 30.71 13.161 ;
 END
 END vss.gds999
 PIN vss.gds1000
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 13.048 33.542 13.248 ;
 END
 END vss.gds1000
 PIN vss.gds1001
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 13.031 31.55 13.231 ;
 END
 END vss.gds1001
 PIN vss.gds1002
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 11.346 33.866 11.546 ;
 END
 END vss.gds1002
 PIN vss.gds1003
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 13.1955 34.886 13.3955 ;
 END
 END vss.gds1003
 PIN vss.gds1004
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 13.1495 34.046 13.3495 ;
 END
 END vss.gds1004
 PIN vss.gds1005
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 10.877 34.366 11.077 ;
 END
 END vss.gds1005
 PIN vss.gds1006
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 31.304 14.679 31.36 14.861 ;
 RECT 32.144 14.739 32.2 14.939 ;
 RECT 31.808 14.698 31.864 14.898 ;
 RECT 31.556 14.679 31.612 14.861 ;
 RECT 32.48 14.698 32.536 14.898 ;
 RECT 33.068 14.698 33.124 14.898 ;
 RECT 32.9 14.698 32.956 14.898 ;
 RECT 33.572 14.679 33.628 14.861 ;
 RECT 33.32 14.679 33.376 14.861 ;
 RECT 34.16 14.698 34.216 14.898 ;
 RECT 34.328 14.698 34.384 14.898 ;
 RECT 30.548 13.354 30.604 13.554 ;
 RECT 31.388 13.354 31.444 13.554 ;
 RECT 30.968 13.354 31.024 13.554 ;
 RECT 31.724 13.335 31.78 13.517 ;
 RECT 31.892 13.354 31.948 13.554 ;
 RECT 33.152 13.335 33.208 13.513 ;
 RECT 32.564 13.354 32.62 13.554 ;
 RECT 32.9 13.335 32.956 13.513 ;
 RECT 33.656 13.354 33.712 13.554 ;
 RECT 34.16 13.354 34.216 13.554 ;
 RECT 34.58 13.354 34.636 13.554 ;
 RECT 30.548 13.074 30.604 13.274 ;
 RECT 30.968 13.074 31.024 13.274 ;
 RECT 31.388 13.074 31.444 13.274 ;
 RECT 31.892 13.074 31.948 13.274 ;
 RECT 31.724 13.111 31.78 13.293 ;
 RECT 32.228 13.0035 32.284 13.2035 ;
 RECT 33.152 13.115 33.208 13.287 ;
 RECT 32.9 13.115 32.956 13.287 ;
 RECT 32.564 13.074 32.62 13.274 ;
 RECT 33.572 13.074 33.628 13.274 ;
 RECT 34.58 13.074 34.636 13.274 ;
 RECT 34.076 13.074 34.132 13.274 ;
 RECT 30.632 10.668 30.688 10.868 ;
 RECT 30.968 10.668 31.024 10.868 ;
 RECT 31.304 10.668 31.36 10.868 ;
 RECT 31.64 10.668 31.696 10.868 ;
 RECT 31.976 10.668 32.032 10.868 ;
 RECT 32.984 10.668 33.04 10.868 ;
 RECT 33.32 10.668 33.376 10.868 ;
 RECT 33.656 10.668 33.712 10.868 ;
 RECT 33.992 10.668 34.048 10.868 ;
 RECT 30.296 11.991 30.352 12.173 ;
 RECT 32.984 12.01 33.04 12.21 ;
 RECT 32.816 12.01 32.872 12.21 ;
 RECT 32.648 12.01 32.704 12.21 ;
 RECT 32.48 12.01 32.536 12.21 ;
 RECT 33.656 12.01 33.712 12.21 ;
 RECT 33.236 11.992 33.292 12.169 ;
 RECT 30.296 11.767 30.352 11.949 ;
 RECT 30.968 11.87 31.024 12.07 ;
 RECT 32.984 11.73 33.04 11.93 ;
 RECT 32.816 11.73 32.872 11.93 ;
 RECT 32.648 11.73 32.704 11.93 ;
 RECT 32.48 11.73 32.536 11.93 ;
 RECT 33.236 11.771 33.292 11.949 ;
 RECT 33.404 11.767 33.46 11.967 ;
 RECT 33.74 11.73 33.796 11.93 ;
 RECT 34.916 11.73 34.972 11.93 ;
 RECT 34.16 11.87 34.216 12.07 ;
 RECT 33.992 11.87 34.048 12.07 ;
 RECT 34.328 11.87 34.384 12.07 ;
 RECT 30.296 10.629 30.352 10.829 ;
 RECT 30.38 13.4245 30.436 13.6245 ;
 RECT 31.22 13.4245 31.276 13.6245 ;
 RECT 30.8 13.4245 30.856 13.6245 ;
 RECT 32.228 13.4245 32.284 13.6245 ;
 RECT 34.832 14.7685 34.888 14.9685 ;
 RECT 34.58 11.9815 34.636 12.1815 ;
 RECT 34.832 12.051 34.888 12.251 ;
 RECT 30.296 14.558 30.352 14.758 ;
 RECT 31.304 14.455 31.36 14.637 ;
 RECT 30.968 14.558 31.024 14.758 ;
 RECT 32.144 14.418 32.2 14.618 ;
 RECT 31.808 14.418 31.864 14.618 ;
 RECT 31.64 14.455 31.696 14.637 ;
 RECT 33.152 14.455 33.208 14.637 ;
 RECT 32.48 14.418 32.536 14.618 ;
 RECT 32.816 14.455 32.872 14.637 ;
 RECT 33.656 14.418 33.712 14.618 ;
 RECT 34.244 14.455 34.3 14.637 ;
 RECT 34.328 10.629 34.384 10.829 ;
 RECT 30.38 10.474 30.436 10.674 ;
 RECT 34.916 10.526 34.972 10.726 ;
 RECT 34.748 10.474 34.804 10.674 ;
 RECT 34.58 10.474 34.636 10.674 ;
 RECT 34.412 10.526 34.468 10.726 ;
 RECT 34.244 10.474 34.3 10.674 ;
 RECT 35.084 10.474 35.14 10.674 ;
 END
 END vss.gds1006
 PIN vss.gds1007
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.102 12.41 40.148 12.61 ;
 END
 END vss.gds1007
 PIN vss.gds1008
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.43 12.41 39.476 12.61 ;
 END
 END vss.gds1008
 PIN vss.gds1009
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.758 12.41 38.804 12.61 ;
 END
 END vss.gds1009
 PIN vss.gds1010
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.086 12.41 38.132 12.61 ;
 END
 END vss.gds1010
 PIN vss.gds1011
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.414 12.41 37.46 12.61 ;
 END
 END vss.gds1011
 PIN vss.gds1012
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.742 12.41 36.788 12.61 ;
 END
 END vss.gds1012
 PIN vss.gds1013
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.07 12.41 36.116 12.61 ;
 END
 END vss.gds1013
 PIN vss.gds1014
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.398 12.41 35.444 12.61 ;
 END
 END vss.gds1014
 PIN vss.gds1015
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.794 12.5875 35.834 12.7875 ;
 END
 END vss.gds1015
 PIN vss.gds1016
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.634 12.105 39.674 12.305 ;
 END
 END vss.gds1016
 PIN vss.gds1017
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.826 12.5875 39.866 12.7875 ;
 END
 END vss.gds1017
 PIN vss.gds1018
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.962 12.105 39.002 12.305 ;
 END
 END vss.gds1018
 PIN vss.gds1019
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.154 12.5875 39.194 12.7875 ;
 END
 END vss.gds1019
 PIN vss.gds1020
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.29 12.105 38.33 12.305 ;
 END
 END vss.gds1020
 PIN vss.gds1021
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.482 12.5875 38.522 12.7875 ;
 END
 END vss.gds1021
 PIN vss.gds1022
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.618 12.105 37.658 12.305 ;
 END
 END vss.gds1022
 PIN vss.gds1023
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 13.1145 37.998 13.3145 ;
 END
 END vss.gds1023
 PIN vss.gds1024
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 13.1145 37.326 13.3145 ;
 END
 END vss.gds1024
 PIN vss.gds1025
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.81 12.5875 37.85 12.7875 ;
 END
 END vss.gds1025
 PIN vss.gds1026
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.946 12.105 36.986 12.305 ;
 END
 END vss.gds1026
 PIN vss.gds1027
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.138 12.5875 37.178 12.7875 ;
 END
 END vss.gds1027
 PIN vss.gds1028
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.274 12.105 36.314 12.305 ;
 END
 END vss.gds1028
 PIN vss.gds1029
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.466 12.5875 36.506 12.7875 ;
 END
 END vss.gds1029
 PIN vss.gds1030
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.602 12.105 35.642 12.305 ;
 END
 END vss.gds1030
 PIN vss.gds1031
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 13.1145 38.67 13.3145 ;
 END
 END vss.gds1031
 PIN vss.gds1032
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 13.1145 36.654 13.3145 ;
 END
 END vss.gds1032
 PIN vss.gds1033
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 13.1145 39.342 13.3145 ;
 END
 END vss.gds1033
 PIN vss.gds1034
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 13.1145 40.014 13.3145 ;
 END
 END vss.gds1034
 PIN vss.gds1035
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 13.1145 35.31 13.3145 ;
 END
 END vss.gds1035
 PIN vss.gds1036
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 13.1145 35.982 13.3145 ;
 END
 END vss.gds1036
 PIN vss.gds1037
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 40.124 12.6525 40.18 12.8525 ;
 RECT 39.62 12.6525 39.676 12.8525 ;
 RECT 39.452 12.6525 39.508 12.8525 ;
 RECT 39.956 12.6525 40.012 12.8525 ;
 RECT 39.788 12.6525 39.844 12.8525 ;
 RECT 38.948 12.6525 39.004 12.8525 ;
 RECT 38.78 12.6525 38.836 12.8525 ;
 RECT 39.284 12.6525 39.34 12.8525 ;
 RECT 39.116 12.6525 39.172 12.8525 ;
 RECT 38.276 12.6525 38.332 12.8525 ;
 RECT 38.108 12.6525 38.164 12.8525 ;
 RECT 38.612 12.6525 38.668 12.8525 ;
 RECT 38.444 12.6525 38.5 12.8525 ;
 RECT 37.604 12.6525 37.66 12.8525 ;
 RECT 37.436 12.6525 37.492 12.8525 ;
 RECT 37.94 12.6525 37.996 12.8525 ;
 RECT 37.772 12.6525 37.828 12.8525 ;
 RECT 36.932 12.6525 36.988 12.8525 ;
 RECT 36.764 12.6525 36.82 12.8525 ;
 RECT 37.268 12.6525 37.324 12.8525 ;
 RECT 37.1 12.6525 37.156 12.8525 ;
 RECT 36.26 12.6525 36.316 12.8525 ;
 RECT 36.092 12.6525 36.148 12.8525 ;
 RECT 36.596 12.6525 36.652 12.8525 ;
 RECT 36.428 12.6525 36.484 12.8525 ;
 RECT 35.588 12.6525 35.644 12.8525 ;
 RECT 35.252 12.6525 35.308 12.8525 ;
 RECT 35.42 12.6525 35.476 12.8525 ;
 RECT 35.924 12.6525 35.98 12.8525 ;
 RECT 35.756 12.6525 35.812 12.8525 ;
 RECT 39.956 14.4275 40.012 14.6275 ;
 RECT 39.284 14.4275 39.34 14.6275 ;
 RECT 38.612 14.4275 38.668 14.6275 ;
 RECT 37.94 14.4275 37.996 14.6275 ;
 RECT 37.268 14.4275 37.324 14.6275 ;
 RECT 36.596 14.4275 36.652 14.6275 ;
 RECT 35.252 14.222 35.308 14.422 ;
 RECT 35.924 14.4275 35.98 14.6275 ;
 RECT 40.124 11.11 40.18 11.31 ;
 RECT 39.62 11.11 39.676 11.31 ;
 RECT 39.452 11.11 39.508 11.31 ;
 RECT 39.788 11.11 39.844 11.31 ;
 RECT 39.956 11.101 40.012 11.301 ;
 RECT 38.948 11.11 39.004 11.31 ;
 RECT 38.78 11.11 38.836 11.31 ;
 RECT 39.116 11.11 39.172 11.31 ;
 RECT 39.284 11.101 39.34 11.301 ;
 RECT 38.276 11.11 38.332 11.31 ;
 RECT 38.108 11.11 38.164 11.31 ;
 RECT 38.444 11.11 38.5 11.31 ;
 RECT 38.612 11.101 38.668 11.301 ;
 RECT 37.604 11.11 37.66 11.31 ;
 RECT 37.436 11.11 37.492 11.31 ;
 RECT 37.772 11.11 37.828 11.31 ;
 RECT 37.94 11.101 37.996 11.301 ;
 RECT 36.932 11.11 36.988 11.31 ;
 RECT 36.764 11.11 36.82 11.31 ;
 RECT 37.1 11.11 37.156 11.31 ;
 RECT 37.268 11.101 37.324 11.301 ;
 RECT 36.26 11.11 36.316 11.31 ;
 RECT 36.092 11.11 36.148 11.31 ;
 RECT 36.428 11.11 36.484 11.31 ;
 RECT 36.596 11.101 36.652 11.301 ;
 RECT 35.252 11.101 35.308 11.301 ;
 RECT 35.588 11.11 35.644 11.31 ;
 RECT 35.42 11.11 35.476 11.31 ;
 RECT 35.756 11.11 35.812 11.31 ;
 RECT 35.924 11.101 35.98 11.301 ;
 END
 END vss.gds1037
 PIN vss.gds1038
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.226 12.41 45.272 12.61 ;
 END
 END vss.gds1038
 PIN vss.gds1039
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.554 12.41 44.6 12.61 ;
 END
 END vss.gds1039
 PIN vss.gds1040
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.882 12.41 43.928 12.61 ;
 END
 END vss.gds1040
 PIN vss.gds1041
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.21 12.41 43.256 12.61 ;
 END
 END vss.gds1041
 PIN vss.gds1042
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.538 12.41 42.584 12.61 ;
 END
 END vss.gds1042
 PIN vss.gds1043
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.866 12.41 41.912 12.61 ;
 END
 END vss.gds1043
 PIN vss.gds1044
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.194 12.41 41.24 12.61 ;
 END
 END vss.gds1044
 PIN vss.gds1045
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.774 13.852 40.814 14.052 ;
 END
 END vss.gds1045
 PIN vss.gds1046
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.918 13.852 40.958 14.052 ;
 END
 END vss.gds1046
 PIN vss.gds1047
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.758 12.105 44.798 12.305 ;
 END
 END vss.gds1047
 PIN vss.gds1048
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.95 12.5875 44.99 12.7875 ;
 END
 END vss.gds1048
 PIN vss.gds1049
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.086 12.105 44.126 12.305 ;
 END
 END vss.gds1049
 PIN vss.gds1050
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.278 12.5875 44.318 12.7875 ;
 END
 END vss.gds1050
 PIN vss.gds1051
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.414 12.105 43.454 12.305 ;
 END
 END vss.gds1051
 PIN vss.gds1052
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.606 12.5875 43.646 12.7875 ;
 END
 END vss.gds1052
 PIN vss.gds1053
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.742 12.105 42.782 12.305 ;
 END
 END vss.gds1053
 PIN vss.gds1054
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.934 12.5875 42.974 12.7875 ;
 END
 END vss.gds1054
 PIN vss.gds1055
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.07 12.105 42.11 12.305 ;
 END
 END vss.gds1055
 PIN vss.gds1056
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.262 12.5875 42.302 12.7875 ;
 END
 END vss.gds1056
 PIN vss.gds1057
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.398 12.105 41.438 12.305 ;
 END
 END vss.gds1057
 PIN vss.gds1058
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.59 12.5875 41.63 12.7875 ;
 END
 END vss.gds1058
 PIN vss.gds1059
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.306 12.105 40.346 12.305 ;
 END
 END vss.gds1059
 PIN vss.gds1060
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.498 12.5875 40.538 12.7875 ;
 END
 END vss.gds1060
 PIN vss.gds1061
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 13.1145 45.138 13.3145 ;
 END
 END vss.gds1061
 PIN vss.gds1062
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 13.1145 44.466 13.3145 ;
 END
 END vss.gds1062
 PIN vss.gds1063
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 13.1145 43.794 13.3145 ;
 END
 END vss.gds1063
 PIN vss.gds1064
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 13.1145 43.122 13.3145 ;
 END
 END vss.gds1064
 PIN vss.gds1065
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 13.1145 42.45 13.3145 ;
 END
 END vss.gds1065
 PIN vss.gds1066
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 13.1145 41.778 13.3145 ;
 END
 END vss.gds1066
 PIN vss.gds1067
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 13.1765 40.686 13.3765 ;
 END
 END vss.gds1067
 PIN vss.gds1068
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.046 13.1765 41.106 13.3765 ;
 END
 END vss.gds1068
 PIN vss.gds1069
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 44.744 12.6525 44.8 12.8525 ;
 RECT 44.576 12.6525 44.632 12.8525 ;
 RECT 45.08 12.6525 45.136 12.8525 ;
 RECT 44.912 12.6525 44.968 12.8525 ;
 RECT 44.072 12.6525 44.128 12.8525 ;
 RECT 43.904 12.6525 43.96 12.8525 ;
 RECT 44.408 12.6525 44.464 12.8525 ;
 RECT 44.24 12.6525 44.296 12.8525 ;
 RECT 43.4 12.6525 43.456 12.8525 ;
 RECT 43.232 12.6525 43.288 12.8525 ;
 RECT 43.736 12.6525 43.792 12.8525 ;
 RECT 43.568 12.6525 43.624 12.8525 ;
 RECT 42.728 12.6525 42.784 12.8525 ;
 RECT 42.56 12.6525 42.616 12.8525 ;
 RECT 43.064 12.6525 43.12 12.8525 ;
 RECT 42.896 12.6525 42.952 12.8525 ;
 RECT 42.056 12.6525 42.112 12.8525 ;
 RECT 41.888 12.6525 41.944 12.8525 ;
 RECT 42.392 12.6525 42.448 12.8525 ;
 RECT 42.224 12.6525 42.28 12.8525 ;
 RECT 41.384 12.6525 41.44 12.8525 ;
 RECT 41.048 12.6525 41.104 12.8525 ;
 RECT 41.216 12.6525 41.272 12.8525 ;
 RECT 41.72 12.6525 41.776 12.8525 ;
 RECT 41.552 12.6525 41.608 12.8525 ;
 RECT 40.628 12.6525 40.684 12.8525 ;
 RECT 40.46 12.6525 40.516 12.8525 ;
 RECT 40.292 12.6525 40.348 12.8525 ;
 RECT 45.08 14.4275 45.136 14.6275 ;
 RECT 44.408 14.4275 44.464 14.6275 ;
 RECT 43.736 14.4275 43.792 14.6275 ;
 RECT 43.064 14.4275 43.12 14.6275 ;
 RECT 42.392 14.4275 42.448 14.6275 ;
 RECT 41.048 14.222 41.104 14.422 ;
 RECT 41.72 14.4275 41.776 14.6275 ;
 RECT 40.628 14.4275 40.684 14.6275 ;
 RECT 44.744 11.11 44.8 11.31 ;
 RECT 44.576 11.11 44.632 11.31 ;
 RECT 44.912 11.11 44.968 11.31 ;
 RECT 45.08 11.101 45.136 11.301 ;
 RECT 44.072 11.11 44.128 11.31 ;
 RECT 43.904 11.11 43.96 11.31 ;
 RECT 44.24 11.11 44.296 11.31 ;
 RECT 44.408 11.101 44.464 11.301 ;
 RECT 43.4 11.11 43.456 11.31 ;
 RECT 43.232 11.11 43.288 11.31 ;
 RECT 43.568 11.11 43.624 11.31 ;
 RECT 43.736 11.101 43.792 11.301 ;
 RECT 42.728 11.11 42.784 11.31 ;
 RECT 42.56 11.11 42.616 11.31 ;
 RECT 42.896 11.11 42.952 11.31 ;
 RECT 43.064 11.101 43.12 11.301 ;
 RECT 42.056 11.11 42.112 11.31 ;
 RECT 41.888 11.11 41.944 11.31 ;
 RECT 42.224 11.11 42.28 11.31 ;
 RECT 42.392 11.101 42.448 11.301 ;
 RECT 41.72 11.101 41.776 11.301 ;
 RECT 40.628 11.101 40.684 11.301 ;
 RECT 41.048 10.9305 41.104 11.1305 ;
 RECT 41.384 11.11 41.44 11.31 ;
 RECT 41.216 11.11 41.272 11.31 ;
 RECT 41.552 11.11 41.608 11.31 ;
 RECT 40.46 11.11 40.516 11.31 ;
 RECT 40.292 11.11 40.348 11.31 ;
 RECT 40.796 12.812 40.852 13.012 ;
 END
 END vss.gds1069
 PIN vss.gds1070
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.898 12.41 45.944 12.61 ;
 END
 END vss.gds1070
 PIN vss.gds1071
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 13.1445 50.25 13.3445 ;
 END
 END vss.gds1071
 PIN vss.gds1072
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.102 12.105 46.142 12.305 ;
 END
 END vss.gds1072
 PIN vss.gds1073
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.294 12.5875 46.334 12.7875 ;
 END
 END vss.gds1073
 PIN vss.gds1074
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.43 12.105 45.47 12.305 ;
 END
 END vss.gds1074
 PIN vss.gds1075
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.622 12.5875 45.662 12.7875 ;
 END
 END vss.gds1075
 PIN vss.gds1076
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 13.1145 45.81 13.3145 ;
 END
 END vss.gds1076
 PIN vss.gds1077
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 12.9745 46.482 13.1745 ;
 END
 END vss.gds1077
 PIN vss.gds1078
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 11.8645 47.162 12.0645 ;
 END
 END vss.gds1078
 PIN vss.gds1079
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.526 11.5435 47.582 11.7435 ;
 END
 END vss.gds1079
 PIN vss.gds1080
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 12.961 46.922 13.161 ;
 END
 END vss.gds1080
 PIN vss.gds1081
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 13.406 46.694 13.606 ;
 END
 END vss.gds1081
 PIN vss.gds1082
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 12.961 47.762 13.161 ;
 END
 END vss.gds1082
 PIN vss.gds1083
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.366 11.488 48.422 11.688 ;
 END
 END vss.gds1083
 PIN vss.gds1084
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 11.699 48.974 11.899 ;
 END
 END vss.gds1084
 PIN vss.gds1085
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 13.0485 49.266 13.2485 ;
 END
 END vss.gds1085
 PIN vss.gds1086
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 13.031 48.602 13.231 ;
 END
 END vss.gds1086
 PIN vss.gds1087
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 13.347 49.946 13.547 ;
 END
 END vss.gds1087
 PIN vss.gds1088
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 11.488 49.522 11.688 ;
 END
 END vss.gds1088
 PIN vss.gds1089
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 46.844 14.698 46.9 14.898 ;
 RECT 48.356 14.679 48.412 14.861 ;
 RECT 49.196 14.739 49.252 14.939 ;
 RECT 48.86 14.698 48.916 14.898 ;
 RECT 48.608 14.679 48.664 14.861 ;
 RECT 49.532 14.698 49.588 14.898 ;
 RECT 50.12 14.698 50.176 14.898 ;
 RECT 49.952 14.698 50.008 14.898 ;
 RECT 47.6 13.354 47.656 13.554 ;
 RECT 48.44 13.354 48.496 13.554 ;
 RECT 48.02 13.354 48.076 13.554 ;
 RECT 48.776 13.335 48.832 13.517 ;
 RECT 48.944 13.354 49 13.554 ;
 RECT 50.204 13.335 50.26 13.513 ;
 RECT 49.616 13.354 49.672 13.554 ;
 RECT 49.952 13.335 50.008 13.513 ;
 RECT 47.6 13.074 47.656 13.274 ;
 RECT 47.18 13.074 47.236 13.274 ;
 RECT 48.02 13.074 48.076 13.274 ;
 RECT 48.44 13.074 48.496 13.274 ;
 RECT 48.944 13.074 49 13.274 ;
 RECT 48.776 13.111 48.832 13.293 ;
 RECT 49.28 13.0035 49.336 13.2035 ;
 RECT 50.204 13.115 50.26 13.287 ;
 RECT 49.952 13.115 50.008 13.287 ;
 RECT 49.616 13.074 49.672 13.274 ;
 RECT 47.684 10.668 47.74 10.868 ;
 RECT 47.012 10.668 47.068 10.868 ;
 RECT 48.02 10.668 48.076 10.868 ;
 RECT 48.356 10.668 48.412 10.868 ;
 RECT 48.692 10.668 48.748 10.868 ;
 RECT 49.028 10.668 49.084 10.868 ;
 RECT 50.036 10.668 50.092 10.868 ;
 RECT 46.76 12.01 46.816 12.21 ;
 RECT 47.348 11.991 47.404 12.173 ;
 RECT 50.036 12.01 50.092 12.21 ;
 RECT 49.868 12.01 49.924 12.21 ;
 RECT 49.7 12.01 49.756 12.21 ;
 RECT 49.532 12.01 49.588 12.21 ;
 RECT 46.76 11.73 46.816 11.93 ;
 RECT 47.348 11.767 47.404 11.949 ;
 RECT 48.02 11.87 48.076 12.07 ;
 RECT 50.036 11.73 50.092 11.93 ;
 RECT 49.868 11.73 49.924 11.93 ;
 RECT 49.7 11.73 49.756 11.93 ;
 RECT 49.532 11.73 49.588 11.93 ;
 RECT 47.348 10.629 47.404 10.829 ;
 RECT 47.18 13.4245 47.236 13.6245 ;
 RECT 47.432 13.4245 47.488 13.6245 ;
 RECT 48.272 13.4245 48.328 13.6245 ;
 RECT 47.852 13.4245 47.908 13.6245 ;
 RECT 49.28 13.4245 49.336 13.6245 ;
 RECT 46.088 12.6525 46.144 12.8525 ;
 RECT 45.92 12.6525 45.976 12.8525 ;
 RECT 46.424 12.6525 46.48 12.8525 ;
 RECT 46.256 12.6525 46.312 12.8525 ;
 RECT 45.416 12.6525 45.472 12.8525 ;
 RECT 45.248 12.6525 45.304 12.8525 ;
 RECT 45.752 12.6525 45.808 12.8525 ;
 RECT 45.584 12.6525 45.64 12.8525 ;
 RECT 47.348 14.558 47.404 14.758 ;
 RECT 48.356 14.455 48.412 14.637 ;
 RECT 48.02 14.558 48.076 14.758 ;
 RECT 49.196 14.418 49.252 14.618 ;
 RECT 48.86 14.418 48.916 14.618 ;
 RECT 48.692 14.455 48.748 14.637 ;
 RECT 50.204 14.455 50.26 14.637 ;
 RECT 49.532 14.418 49.588 14.618 ;
 RECT 49.868 14.455 49.924 14.637 ;
 RECT 46.424 14.4275 46.48 14.6275 ;
 RECT 45.752 14.4275 45.808 14.6275 ;
 RECT 46.088 11.11 46.144 11.31 ;
 RECT 46.424 11.101 46.48 11.301 ;
 RECT 45.416 11.11 45.472 11.31 ;
 RECT 45.248 11.11 45.304 11.31 ;
 RECT 45.584 11.11 45.64 11.31 ;
 RECT 45.752 11.101 45.808 11.301 ;
 RECT 45.92 11.11 45.976 11.31 ;
 RECT 46.256 11.11 46.312 11.31 ;
 RECT 47.432 10.474 47.488 10.674 ;
 RECT 47.264 10.474 47.32 10.674 ;
 RECT 46.928 10.474 46.984 10.674 ;
 RECT 46.592 10.474 46.648 10.674 ;
 RECT 47.096 10.474 47.152 10.674 ;
 RECT 46.76 10.5945 46.816 10.7945 ;
 END
 END vss.gds1089
 PIN vss.gds1090
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.138 12.41 55.184 12.61 ;
 END
 END vss.gds1090
 PIN vss.gds1091
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.466 12.41 54.512 12.61 ;
 END
 END vss.gds1091
 PIN vss.gds1092
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.794 12.41 53.84 12.61 ;
 END
 END vss.gds1092
 PIN vss.gds1093
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.122 12.41 53.168 12.61 ;
 END
 END vss.gds1093
 PIN vss.gds1094
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.45 12.41 52.496 12.61 ;
 END
 END vss.gds1094
 PIN vss.gds1095
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.698 14.951 50.754 15.151 ;
 END
 END vss.gds1095
 PIN vss.gds1096
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.846 12.5875 52.886 12.7875 ;
 END
 END vss.gds1096
 PIN vss.gds1097
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 14.29 51.418 14.49 ;
 END
 END vss.gds1097
 PIN vss.gds1098
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.702 13.515 51.758 13.715 ;
 END
 END vss.gds1098
 PIN vss.gds1099
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.67 12.105 54.71 12.305 ;
 END
 END vss.gds1099
 PIN vss.gds1100
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.862 12.5875 54.902 12.7875 ;
 END
 END vss.gds1100
 PIN vss.gds1101
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.998 12.105 54.038 12.305 ;
 END
 END vss.gds1101
 PIN vss.gds1102
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 13.1145 54.378 13.3145 ;
 END
 END vss.gds1102
 PIN vss.gds1103
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 13.1145 55.05 13.3145 ;
 END
 END vss.gds1103
 PIN vss.gds1104
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 13.1145 53.706 13.3145 ;
 END
 END vss.gds1104
 PIN vss.gds1105
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.19 12.5875 54.23 12.7875 ;
 END
 END vss.gds1105
 PIN vss.gds1106
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.326 12.105 53.366 12.305 ;
 END
 END vss.gds1106
 PIN vss.gds1107
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.518 12.5875 53.558 12.7875 ;
 END
 END vss.gds1107
 PIN vss.gds1108
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.654 12.105 52.694 12.305 ;
 END
 END vss.gds1108
 PIN vss.gds1109
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 10.877 51.418 11.077 ;
 END
 END vss.gds1109
 PIN vss.gds1110
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.274 14.5535 50.33 14.7535 ;
 END
 END vss.gds1110
 PIN vss.gds1111
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 11.346 50.918 11.546 ;
 END
 END vss.gds1111
 PIN vss.gds1112
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 13.1145 53.034 13.3145 ;
 END
 END vss.gds1112
 PIN vss.gds1113
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 13.1955 51.938 13.3955 ;
 END
 END vss.gds1113
 PIN vss.gds1114
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 13.048 50.594 13.248 ;
 END
 END vss.gds1114
 PIN vss.gds1115
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 13.1145 52.362 13.3145 ;
 END
 END vss.gds1115
 PIN vss.gds1116
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 13.1495 51.098 13.3495 ;
 END
 END vss.gds1116
 PIN vss.gds1117
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 50.624 14.679 50.68 14.861 ;
 RECT 50.372 14.679 50.428 14.861 ;
 RECT 51.212 14.698 51.268 14.898 ;
 RECT 51.38 14.698 51.436 14.898 ;
 RECT 50.708 13.354 50.764 13.554 ;
 RECT 51.212 13.354 51.268 13.554 ;
 RECT 51.632 13.354 51.688 13.554 ;
 RECT 50.624 13.074 50.68 13.274 ;
 RECT 51.632 13.074 51.688 13.274 ;
 RECT 51.128 13.074 51.184 13.274 ;
 RECT 50.372 10.668 50.428 10.868 ;
 RECT 50.708 10.668 50.764 10.868 ;
 RECT 51.044 10.668 51.1 10.868 ;
 RECT 50.708 12.01 50.764 12.21 ;
 RECT 50.288 11.992 50.344 12.169 ;
 RECT 50.288 11.771 50.344 11.949 ;
 RECT 50.456 11.767 50.512 11.967 ;
 RECT 50.792 11.73 50.848 11.93 ;
 RECT 51.968 11.73 52.024 11.93 ;
 RECT 52.304 14.222 52.36 14.422 ;
 RECT 51.212 11.87 51.268 12.07 ;
 RECT 51.044 11.87 51.1 12.07 ;
 RECT 51.38 11.87 51.436 12.07 ;
 RECT 55.16 12.6525 55.216 12.8525 ;
 RECT 54.656 12.6525 54.712 12.8525 ;
 RECT 54.488 12.6525 54.544 12.8525 ;
 RECT 54.992 12.6525 55.048 12.8525 ;
 RECT 54.824 12.6525 54.88 12.8525 ;
 RECT 53.984 12.6525 54.04 12.8525 ;
 RECT 53.816 12.6525 53.872 12.8525 ;
 RECT 54.32 12.6525 54.376 12.8525 ;
 RECT 54.152 12.6525 54.208 12.8525 ;
 RECT 53.312 12.6525 53.368 12.8525 ;
 RECT 53.144 12.6525 53.2 12.8525 ;
 RECT 53.648 12.6525 53.704 12.8525 ;
 RECT 53.48 12.6525 53.536 12.8525 ;
 RECT 52.64 12.6525 52.696 12.8525 ;
 RECT 52.304 12.6525 52.36 12.8525 ;
 RECT 52.472 12.6525 52.528 12.8525 ;
 RECT 52.976 12.6525 53.032 12.8525 ;
 RECT 52.808 12.6525 52.864 12.8525 ;
 RECT 51.884 14.7685 51.94 14.9685 ;
 RECT 51.632 11.9815 51.688 12.1815 ;
 RECT 51.884 12.051 51.94 12.251 ;
 RECT 54.992 14.4275 55.048 14.6275 ;
 RECT 54.32 14.4275 54.376 14.6275 ;
 RECT 53.648 14.4275 53.704 14.6275 ;
 RECT 52.976 14.4275 53.032 14.6275 ;
 RECT 50.708 14.418 50.764 14.618 ;
 RECT 51.296 14.455 51.352 14.637 ;
 RECT 55.16 11.11 55.216 11.31 ;
 RECT 54.656 11.11 54.712 11.31 ;
 RECT 54.488 11.11 54.544 11.31 ;
 RECT 54.824 11.11 54.88 11.31 ;
 RECT 54.992 11.101 55.048 11.301 ;
 RECT 53.984 11.11 54.04 11.31 ;
 RECT 53.816 11.11 53.872 11.31 ;
 RECT 54.152 11.11 54.208 11.31 ;
 RECT 54.32 11.101 54.376 11.301 ;
 RECT 53.312 11.11 53.368 11.31 ;
 RECT 53.144 11.11 53.2 11.31 ;
 RECT 53.48 11.11 53.536 11.31 ;
 RECT 53.648 11.101 53.704 11.301 ;
 RECT 52.304 11.101 52.36 11.301 ;
 RECT 51.38 10.629 51.436 10.829 ;
 RECT 52.64 11.11 52.696 11.31 ;
 RECT 52.472 11.11 52.528 11.31 ;
 RECT 52.808 11.11 52.864 11.31 ;
 RECT 52.976 11.101 53.032 11.301 ;
 RECT 51.968 10.526 52.024 10.726 ;
 RECT 51.8 10.474 51.856 10.674 ;
 RECT 51.632 10.474 51.688 10.674 ;
 RECT 51.464 10.526 51.52 10.726 ;
 RECT 51.296 10.474 51.352 10.674 ;
 RECT 52.136 10.474 52.192 10.674 ;
 END
 END vss.gds1117
 PIN vss.gds1118
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.59 12.41 59.636 12.61 ;
 END
 END vss.gds1118
 PIN vss.gds1119
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.918 12.41 58.964 12.61 ;
 END
 END vss.gds1119
 PIN vss.gds1120
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.246 12.41 58.292 12.61 ;
 END
 END vss.gds1120
 PIN vss.gds1121
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.154 12.41 57.2 12.61 ;
 END
 END vss.gds1121
 PIN vss.gds1122
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.482 12.41 56.528 12.61 ;
 END
 END vss.gds1122
 PIN vss.gds1123
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.81 12.41 55.856 12.61 ;
 END
 END vss.gds1123
 PIN vss.gds1124
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.826 13.852 57.866 14.052 ;
 END
 END vss.gds1124
 PIN vss.gds1125
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.97 13.852 58.01 14.052 ;
 END
 END vss.gds1125
 PIN vss.gds1126
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.098 13.1765 58.158 13.3765 ;
 END
 END vss.gds1126
 PIN vss.gds1127
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.794 12.105 59.834 12.305 ;
 END
 END vss.gds1127
 PIN vss.gds1128
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.986 12.5875 60.026 12.7875 ;
 END
 END vss.gds1128
 PIN vss.gds1129
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.122 12.105 59.162 12.305 ;
 END
 END vss.gds1129
 PIN vss.gds1130
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.314 12.5875 59.354 12.7875 ;
 END
 END vss.gds1130
 PIN vss.gds1131
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.45 12.105 58.49 12.305 ;
 END
 END vss.gds1131
 PIN vss.gds1132
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.642 12.5875 58.682 12.7875 ;
 END
 END vss.gds1132
 PIN vss.gds1133
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.358 12.105 57.398 12.305 ;
 END
 END vss.gds1133
 PIN vss.gds1134
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.55 12.5875 57.59 12.7875 ;
 END
 END vss.gds1134
 PIN vss.gds1135
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.686 12.105 56.726 12.305 ;
 END
 END vss.gds1135
 PIN vss.gds1136
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.878 12.5875 56.918 12.7875 ;
 END
 END vss.gds1136
 PIN vss.gds1137
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.014 12.105 56.054 12.305 ;
 END
 END vss.gds1137
 PIN vss.gds1138
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.206 12.5875 56.246 12.7875 ;
 END
 END vss.gds1138
 PIN vss.gds1139
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.342 12.105 55.382 12.305 ;
 END
 END vss.gds1139
 PIN vss.gds1140
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.534 12.5875 55.574 12.7875 ;
 END
 END vss.gds1140
 PIN vss.gds1141
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 13.1145 60.174 13.3145 ;
 END
 END vss.gds1141
 PIN vss.gds1142
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 13.1145 59.502 13.3145 ;
 END
 END vss.gds1142
 PIN vss.gds1143
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 13.1145 58.83 13.3145 ;
 END
 END vss.gds1143
 PIN vss.gds1144
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 13.1145 55.722 13.3145 ;
 END
 END vss.gds1144
 PIN vss.gds1145
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 13.1145 56.394 13.3145 ;
 END
 END vss.gds1145
 PIN vss.gds1146
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 13.1765 57.738 13.3765 ;
 END
 END vss.gds1146
 PIN vss.gds1147
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 13.1145 57.066 13.3145 ;
 END
 END vss.gds1147
 PIN vss.gds1148
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 59.78 11.11 59.836 11.31 ;
 RECT 59.612 11.11 59.668 11.31 ;
 RECT 59.948 11.11 60.004 11.31 ;
 RECT 60.116 11.101 60.172 11.301 ;
 RECT 59.108 11.11 59.164 11.31 ;
 RECT 58.94 11.11 58.996 11.31 ;
 RECT 59.276 11.11 59.332 11.31 ;
 RECT 59.444 11.101 59.5 11.301 ;
 RECT 58.772 11.101 58.828 11.301 ;
 RECT 58.1 10.9305 58.156 11.1305 ;
 RECT 58.436 11.11 58.492 11.31 ;
 RECT 58.268 11.11 58.324 11.31 ;
 RECT 58.604 11.11 58.66 11.31 ;
 RECT 58.1 14.222 58.156 14.422 ;
 RECT 59.78 12.6525 59.836 12.8525 ;
 RECT 59.612 12.6525 59.668 12.8525 ;
 RECT 60.116 12.6525 60.172 12.8525 ;
 RECT 59.948 12.6525 60.004 12.8525 ;
 RECT 59.108 12.6525 59.164 12.8525 ;
 RECT 58.94 12.6525 58.996 12.8525 ;
 RECT 59.444 12.6525 59.5 12.8525 ;
 RECT 59.276 12.6525 59.332 12.8525 ;
 RECT 58.436 12.6525 58.492 12.8525 ;
 RECT 58.1 12.6525 58.156 12.8525 ;
 RECT 58.268 12.6525 58.324 12.8525 ;
 RECT 58.772 12.6525 58.828 12.8525 ;
 RECT 58.604 12.6525 58.66 12.8525 ;
 RECT 57.344 12.6525 57.4 12.8525 ;
 RECT 57.176 12.6525 57.232 12.8525 ;
 RECT 57.68 12.6525 57.736 12.8525 ;
 RECT 57.512 12.6525 57.568 12.8525 ;
 RECT 56.672 12.6525 56.728 12.8525 ;
 RECT 56.504 12.6525 56.56 12.8525 ;
 RECT 57.008 12.6525 57.064 12.8525 ;
 RECT 56.84 12.6525 56.896 12.8525 ;
 RECT 56 12.6525 56.056 12.8525 ;
 RECT 55.832 12.6525 55.888 12.8525 ;
 RECT 56.336 12.6525 56.392 12.8525 ;
 RECT 56.168 12.6525 56.224 12.8525 ;
 RECT 55.328 12.6525 55.384 12.8525 ;
 RECT 55.664 12.6525 55.72 12.8525 ;
 RECT 55.496 12.6525 55.552 12.8525 ;
 RECT 60.116 14.4275 60.172 14.6275 ;
 RECT 59.444 14.4275 59.5 14.6275 ;
 RECT 58.772 14.4275 58.828 14.6275 ;
 RECT 57.68 14.4275 57.736 14.6275 ;
 RECT 57.008 14.4275 57.064 14.6275 ;
 RECT 56.336 14.4275 56.392 14.6275 ;
 RECT 55.664 14.4275 55.72 14.6275 ;
 RECT 57.344 11.11 57.4 11.31 ;
 RECT 57.176 11.11 57.232 11.31 ;
 RECT 57.512 11.11 57.568 11.31 ;
 RECT 57.68 11.101 57.736 11.301 ;
 RECT 56.672 11.11 56.728 11.31 ;
 RECT 56.504 11.11 56.56 11.31 ;
 RECT 56.84 11.11 56.896 11.31 ;
 RECT 57.008 11.101 57.064 11.301 ;
 RECT 56 11.11 56.056 11.31 ;
 RECT 55.832 11.11 55.888 11.31 ;
 RECT 56.168 11.11 56.224 11.31 ;
 RECT 56.336 11.101 56.392 11.301 ;
 RECT 55.328 11.11 55.384 11.31 ;
 RECT 55.496 11.11 55.552 11.31 ;
 RECT 55.664 11.101 55.72 11.301 ;
 RECT 57.848 12.812 57.904 13.012 ;
 END
 END vss.gds1148
 PIN vss.gds1149
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.95 12.41 62.996 12.61 ;
 END
 END vss.gds1149
 PIN vss.gds1150
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.278 12.41 62.324 12.61 ;
 END
 END vss.gds1150
 PIN vss.gds1151
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.606 12.41 61.652 12.61 ;
 END
 END vss.gds1151
 PIN vss.gds1152
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.934 12.41 60.98 12.61 ;
 END
 END vss.gds1152
 PIN vss.gds1153
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.262 12.41 60.308 12.61 ;
 END
 END vss.gds1153
 PIN vss.gds1154
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 11.8645 64.214 12.0645 ;
 END
 END vss.gds1154
 PIN vss.gds1155
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.578 11.5435 64.634 11.7435 ;
 END
 END vss.gds1155
 PIN vss.gds1156
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.154 12.105 63.194 12.305 ;
 END
 END vss.gds1156
 PIN vss.gds1157
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.346 12.5875 63.386 12.7875 ;
 END
 END vss.gds1157
 PIN vss.gds1158
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.482 12.105 62.522 12.305 ;
 END
 END vss.gds1158
 PIN vss.gds1159
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.674 12.5875 62.714 12.7875 ;
 END
 END vss.gds1159
 PIN vss.gds1160
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.81 12.105 61.85 12.305 ;
 END
 END vss.gds1160
 PIN vss.gds1161
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.002 12.5875 62.042 12.7875 ;
 END
 END vss.gds1161
 PIN vss.gds1162
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.138 12.105 61.178 12.305 ;
 END
 END vss.gds1162
 PIN vss.gds1163
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.33 12.5875 61.37 12.7875 ;
 END
 END vss.gds1163
 PIN vss.gds1164
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.466 12.105 60.506 12.305 ;
 END
 END vss.gds1164
 PIN vss.gds1165
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.658 12.5875 60.698 12.7875 ;
 END
 END vss.gds1165
 PIN vss.gds1166
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 12.9745 63.534 13.1745 ;
 END
 END vss.gds1166
 PIN vss.gds1167
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 13.1145 62.862 13.3145 ;
 END
 END vss.gds1167
 PIN vss.gds1168
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 13.1145 62.19 13.3145 ;
 END
 END vss.gds1168
 PIN vss.gds1169
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 13.1145 61.518 13.3145 ;
 END
 END vss.gds1169
 PIN vss.gds1170
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 13.1145 60.846 13.3145 ;
 END
 END vss.gds1170
 PIN vss.gds1171
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 12.961 63.974 13.161 ;
 END
 END vss.gds1171
 PIN vss.gds1172
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 13.406 63.746 13.606 ;
 END
 END vss.gds1172
 PIN vss.gds1173
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 12.961 64.814 13.161 ;
 END
 END vss.gds1173
 PIN vss.gds1174
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 63.896 14.698 63.952 14.898 ;
 RECT 64.652 13.354 64.708 13.554 ;
 RECT 65.072 13.354 65.128 13.554 ;
 RECT 64.652 13.074 64.708 13.274 ;
 RECT 64.232 13.074 64.288 13.274 ;
 RECT 65.072 13.074 65.128 13.274 ;
 RECT 64.736 10.668 64.792 10.868 ;
 RECT 64.064 10.668 64.12 10.868 ;
 RECT 65.072 10.668 65.128 10.868 ;
 RECT 63.812 12.01 63.868 12.21 ;
 RECT 64.4 11.991 64.456 12.173 ;
 RECT 63.812 11.73 63.868 11.93 ;
 RECT 64.4 11.767 64.456 11.949 ;
 RECT 65.072 11.87 65.128 12.07 ;
 RECT 64.4 10.629 64.456 10.829 ;
 RECT 63.14 11.11 63.196 11.31 ;
 RECT 63.476 11.101 63.532 11.301 ;
 RECT 62.468 11.11 62.524 11.31 ;
 RECT 62.3 11.11 62.356 11.31 ;
 RECT 62.636 11.11 62.692 11.31 ;
 RECT 62.804 11.101 62.86 11.301 ;
 RECT 61.796 11.11 61.852 11.31 ;
 RECT 61.628 11.11 61.684 11.31 ;
 RECT 61.964 11.11 62.02 11.31 ;
 RECT 62.132 11.101 62.188 11.301 ;
 RECT 61.124 11.11 61.18 11.31 ;
 RECT 60.956 11.11 61.012 11.31 ;
 RECT 61.292 11.11 61.348 11.31 ;
 RECT 61.46 11.101 61.516 11.301 ;
 RECT 60.788 11.101 60.844 11.301 ;
 RECT 60.452 11.11 60.508 11.31 ;
 RECT 60.62 11.11 60.676 11.31 ;
 RECT 60.284 11.11 60.34 11.31 ;
 RECT 63.14 12.6525 63.196 12.8525 ;
 RECT 62.972 12.6525 63.028 12.8525 ;
 RECT 63.476 12.6525 63.532 12.8525 ;
 RECT 63.308 12.6525 63.364 12.8525 ;
 RECT 62.468 12.6525 62.524 12.8525 ;
 RECT 62.3 12.6525 62.356 12.8525 ;
 RECT 62.804 12.6525 62.86 12.8525 ;
 RECT 62.636 12.6525 62.692 12.8525 ;
 RECT 61.796 12.6525 61.852 12.8525 ;
 RECT 61.628 12.6525 61.684 12.8525 ;
 RECT 62.132 12.6525 62.188 12.8525 ;
 RECT 61.964 12.6525 62.02 12.8525 ;
 RECT 61.124 12.6525 61.18 12.8525 ;
 RECT 60.956 12.6525 61.012 12.8525 ;
 RECT 61.46 12.6525 61.516 12.8525 ;
 RECT 61.292 12.6525 61.348 12.8525 ;
 RECT 60.452 12.6525 60.508 12.8525 ;
 RECT 60.788 12.6525 60.844 12.8525 ;
 RECT 60.62 12.6525 60.676 12.8525 ;
 RECT 60.284 12.6525 60.34 12.8525 ;
 RECT 64.232 13.4245 64.288 13.6245 ;
 RECT 64.484 13.4245 64.54 13.6245 ;
 RECT 64.904 13.4245 64.96 13.6245 ;
 RECT 63.476 14.4275 63.532 14.6275 ;
 RECT 62.804 14.4275 62.86 14.6275 ;
 RECT 62.132 14.4275 62.188 14.6275 ;
 RECT 61.46 14.4275 61.516 14.6275 ;
 RECT 60.788 14.4275 60.844 14.6275 ;
 RECT 64.4 14.558 64.456 14.758 ;
 RECT 65.072 14.558 65.128 14.758 ;
 RECT 64.484 10.474 64.54 10.674 ;
 RECT 63.98 10.474 64.036 10.674 ;
 RECT 64.316 10.474 64.372 10.674 ;
 RECT 64.148 10.474 64.204 10.674 ;
 RECT 63.644 10.474 63.7 10.674 ;
 RECT 62.972 11.11 63.028 11.31 ;
 RECT 63.308 11.11 63.364 11.31 ;
 RECT 63.812 10.5945 63.868 10.7945 ;
 END
 END vss.gds1174
 PIN vss.gds1175
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.174 12.41 70.22 12.61 ;
 END
 END vss.gds1175
 PIN vss.gds1176
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.502 12.41 69.548 12.61 ;
 END
 END vss.gds1176
 PIN vss.gds1177
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.898 12.5875 69.938 12.7875 ;
 END
 END vss.gds1177
 PIN vss.gds1178
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.75 14.951 67.806 15.151 ;
 END
 END vss.gds1178
 PIN vss.gds1179
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.326 14.5535 67.382 14.7535 ;
 END
 END vss.gds1179
 PIN vss.gds1180
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 13.1445 67.302 13.3445 ;
 END
 END vss.gds1180
 PIN vss.gds1181
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 14.29 68.47 14.49 ;
 END
 END vss.gds1181
 PIN vss.gds1182
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.754 13.515 68.81 13.715 ;
 END
 END vss.gds1182
 PIN vss.gds1183
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.418 11.488 65.474 11.688 ;
 END
 END vss.gds1183
 PIN vss.gds1184
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 11.699 66.026 11.899 ;
 END
 END vss.gds1184
 PIN vss.gds1185
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 11.488 66.574 11.688 ;
 END
 END vss.gds1185
 PIN vss.gds1186
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 13.0485 66.318 13.2485 ;
 END
 END vss.gds1186
 PIN vss.gds1187
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 13.1145 70.086 13.3145 ;
 END
 END vss.gds1187
 PIN vss.gds1188
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 13.1495 68.15 13.3495 ;
 END
 END vss.gds1188
 PIN vss.gds1189
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 13.048 67.646 13.248 ;
 END
 END vss.gds1189
 PIN vss.gds1190
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.706 12.105 69.746 12.305 ;
 END
 END vss.gds1190
 PIN vss.gds1191
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 11.346 67.97 11.546 ;
 END
 END vss.gds1191
 PIN vss.gds1192
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 13.031 65.654 13.231 ;
 END
 END vss.gds1192
 PIN vss.gds1193
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 13.347 66.998 13.547 ;
 END
 END vss.gds1193
 PIN vss.gds1194
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 13.1955 68.99 13.3955 ;
 END
 END vss.gds1194
 PIN vss.gds1195
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 10.877 68.47 11.077 ;
 END
 END vss.gds1195
 PIN vss.gds1196
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 13.1145 69.414 13.3145 ;
 END
 END vss.gds1196
 PIN vss.gds1197
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 65.408 14.679 65.464 14.861 ;
 RECT 66.248 14.739 66.304 14.939 ;
 RECT 65.912 14.698 65.968 14.898 ;
 RECT 65.66 14.679 65.716 14.861 ;
 RECT 66.584 14.698 66.64 14.898 ;
 RECT 67.172 14.698 67.228 14.898 ;
 RECT 67.004 14.698 67.06 14.898 ;
 RECT 67.676 14.679 67.732 14.861 ;
 RECT 67.424 14.679 67.48 14.861 ;
 RECT 68.264 14.698 68.32 14.898 ;
 RECT 68.432 14.698 68.488 14.898 ;
 RECT 65.492 13.354 65.548 13.554 ;
 RECT 65.828 13.335 65.884 13.517 ;
 RECT 65.996 13.354 66.052 13.554 ;
 RECT 67.256 13.335 67.312 13.513 ;
 RECT 66.668 13.354 66.724 13.554 ;
 RECT 67.004 13.335 67.06 13.513 ;
 RECT 67.76 13.354 67.816 13.554 ;
 RECT 68.264 13.354 68.32 13.554 ;
 RECT 68.684 13.354 68.74 13.554 ;
 RECT 65.492 13.074 65.548 13.274 ;
 RECT 65.996 13.074 66.052 13.274 ;
 RECT 65.828 13.111 65.884 13.293 ;
 RECT 66.332 13.0035 66.388 13.2035 ;
 RECT 67.256 13.115 67.312 13.287 ;
 RECT 67.004 13.115 67.06 13.287 ;
 RECT 66.668 13.074 66.724 13.274 ;
 RECT 67.676 13.074 67.732 13.274 ;
 RECT 68.684 13.074 68.74 13.274 ;
 RECT 68.18 13.074 68.236 13.274 ;
 RECT 65.408 10.668 65.464 10.868 ;
 RECT 65.744 10.668 65.8 10.868 ;
 RECT 66.08 10.668 66.136 10.868 ;
 RECT 67.088 10.668 67.144 10.868 ;
 RECT 67.424 10.668 67.48 10.868 ;
 RECT 67.76 10.668 67.816 10.868 ;
 RECT 68.096 10.668 68.152 10.868 ;
 RECT 67.088 12.01 67.144 12.21 ;
 RECT 66.92 12.01 66.976 12.21 ;
 RECT 66.752 12.01 66.808 12.21 ;
 RECT 66.584 12.01 66.64 12.21 ;
 RECT 67.76 12.01 67.816 12.21 ;
 RECT 67.34 11.992 67.396 12.169 ;
 RECT 67.088 11.73 67.144 11.93 ;
 RECT 66.92 11.73 66.976 11.93 ;
 RECT 66.752 11.73 66.808 11.93 ;
 RECT 66.584 11.73 66.64 11.93 ;
 RECT 67.34 11.771 67.396 11.949 ;
 RECT 67.508 11.767 67.564 11.967 ;
 RECT 67.844 11.73 67.9 11.93 ;
 RECT 69.02 11.73 69.076 11.93 ;
 RECT 68.264 11.87 68.32 12.07 ;
 RECT 68.096 11.87 68.152 12.07 ;
 RECT 68.432 11.87 68.488 12.07 ;
 RECT 65.324 13.4245 65.38 13.6245 ;
 RECT 66.332 13.4245 66.388 13.6245 ;
 RECT 70.196 11.11 70.252 11.31 ;
 RECT 69.356 11.101 69.412 11.301 ;
 RECT 68.432 10.629 68.488 10.829 ;
 RECT 69.692 11.11 69.748 11.31 ;
 RECT 69.524 11.11 69.58 11.31 ;
 RECT 69.86 11.11 69.916 11.31 ;
 RECT 70.028 11.101 70.084 11.301 ;
 RECT 68.936 14.7685 68.992 14.9685 ;
 RECT 65.408 14.455 65.464 14.637 ;
 RECT 66.248 14.418 66.304 14.618 ;
 RECT 65.912 14.418 65.968 14.618 ;
 RECT 65.744 14.455 65.8 14.637 ;
 RECT 67.256 14.455 67.312 14.637 ;
 RECT 66.584 14.418 66.64 14.618 ;
 RECT 66.92 14.455 66.976 14.637 ;
 RECT 67.76 14.418 67.816 14.618 ;
 RECT 68.348 14.455 68.404 14.637 ;
 RECT 70.196 12.6525 70.252 12.8525 ;
 RECT 69.692 12.6525 69.748 12.8525 ;
 RECT 69.356 12.6525 69.412 12.8525 ;
 RECT 69.524 12.6525 69.58 12.8525 ;
 RECT 70.028 12.6525 70.084 12.8525 ;
 RECT 69.86 12.6525 69.916 12.8525 ;
 RECT 68.684 11.9815 68.74 12.1815 ;
 RECT 68.936 12.051 68.992 12.251 ;
 RECT 69.356 14.222 69.412 14.422 ;
 RECT 70.028 14.4275 70.084 14.6275 ;
 RECT 69.02 10.526 69.076 10.726 ;
 RECT 68.852 10.474 68.908 10.674 ;
 RECT 68.684 10.474 68.74 10.674 ;
 RECT 68.516 10.526 68.572 10.726 ;
 RECT 68.348 10.474 68.404 10.674 ;
 RECT 69.188 10.474 69.244 10.674 ;
 END
 END vss.gds1197
 PIN vss.gds1198
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.206 12.41 74.252 12.61 ;
 END
 END vss.gds1198
 PIN vss.gds1199
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.534 12.41 73.58 12.61 ;
 END
 END vss.gds1199
 PIN vss.gds1200
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.862 12.41 72.908 12.61 ;
 END
 END vss.gds1200
 PIN vss.gds1201
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.19 12.41 72.236 12.61 ;
 END
 END vss.gds1201
 PIN vss.gds1202
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.518 12.41 71.564 12.61 ;
 END
 END vss.gds1202
 PIN vss.gds1203
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.846 12.41 70.892 12.61 ;
 END
 END vss.gds1203
 PIN vss.gds1204
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.41 12.105 74.45 12.305 ;
 END
 END vss.gds1204
 PIN vss.gds1205
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.602 12.5875 74.642 12.7875 ;
 END
 END vss.gds1205
 PIN vss.gds1206
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.738 12.105 73.778 12.305 ;
 END
 END vss.gds1206
 PIN vss.gds1207
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.93 12.5875 73.97 12.7875 ;
 END
 END vss.gds1207
 PIN vss.gds1208
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.066 12.105 73.106 12.305 ;
 END
 END vss.gds1208
 PIN vss.gds1209
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.258 12.5875 73.298 12.7875 ;
 END
 END vss.gds1209
 PIN vss.gds1210
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.394 12.105 72.434 12.305 ;
 END
 END vss.gds1210
 PIN vss.gds1211
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.586 12.5875 72.626 12.7875 ;
 END
 END vss.gds1211
 PIN vss.gds1212
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.722 12.105 71.762 12.305 ;
 END
 END vss.gds1212
 PIN vss.gds1213
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.914 12.5875 71.954 12.7875 ;
 END
 END vss.gds1213
 PIN vss.gds1214
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.05 12.105 71.09 12.305 ;
 END
 END vss.gds1214
 PIN vss.gds1215
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.242 12.5875 71.282 12.7875 ;
 END
 END vss.gds1215
 PIN vss.gds1216
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 13.1145 71.43 13.3145 ;
 END
 END vss.gds1216
 PIN vss.gds1217
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 13.1145 72.102 13.3145 ;
 END
 END vss.gds1217
 PIN vss.gds1218
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 13.1145 72.774 13.3145 ;
 END
 END vss.gds1218
 PIN vss.gds1219
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 13.1145 70.758 13.3145 ;
 END
 END vss.gds1219
 PIN vss.gds1220
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.378 12.105 70.418 12.305 ;
 END
 END vss.gds1220
 PIN vss.gds1221
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.57 12.5875 70.61 12.7875 ;
 END
 END vss.gds1221
 PIN vss.gds1222
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 13.1145 74.118 13.3145 ;
 END
 END vss.gds1222
 PIN vss.gds1223
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 13.1145 74.79 13.3145 ;
 END
 END vss.gds1223
 PIN vss.gds1224
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 13.1145 73.446 13.3145 ;
 END
 END vss.gds1224
 PIN vss.gds1225
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 74.396 11.11 74.452 11.31 ;
 RECT 74.228 11.11 74.284 11.31 ;
 RECT 74.564 11.11 74.62 11.31 ;
 RECT 74.732 11.101 74.788 11.301 ;
 RECT 73.724 11.11 73.78 11.31 ;
 RECT 73.556 11.11 73.612 11.31 ;
 RECT 73.892 11.11 73.948 11.31 ;
 RECT 74.06 11.101 74.116 11.301 ;
 RECT 73.052 11.11 73.108 11.31 ;
 RECT 72.884 11.11 72.94 11.31 ;
 RECT 73.22 11.11 73.276 11.31 ;
 RECT 73.388 11.101 73.444 11.301 ;
 RECT 72.38 11.11 72.436 11.31 ;
 RECT 72.212 11.11 72.268 11.31 ;
 RECT 72.548 11.11 72.604 11.31 ;
 RECT 72.716 11.101 72.772 11.301 ;
 RECT 71.708 11.11 71.764 11.31 ;
 RECT 71.54 11.11 71.596 11.31 ;
 RECT 71.876 11.11 71.932 11.31 ;
 RECT 72.044 11.101 72.1 11.301 ;
 RECT 71.036 11.11 71.092 11.31 ;
 RECT 70.868 11.11 70.924 11.31 ;
 RECT 71.204 11.11 71.26 11.31 ;
 RECT 71.372 11.101 71.428 11.301 ;
 RECT 70.364 11.11 70.42 11.31 ;
 RECT 70.532 11.11 70.588 11.31 ;
 RECT 70.7 11.101 70.756 11.301 ;
 RECT 74.396 12.6525 74.452 12.8525 ;
 RECT 74.228 12.6525 74.284 12.8525 ;
 RECT 74.732 12.6525 74.788 12.8525 ;
 RECT 74.564 12.6525 74.62 12.8525 ;
 RECT 73.724 12.6525 73.78 12.8525 ;
 RECT 73.556 12.6525 73.612 12.8525 ;
 RECT 74.06 12.6525 74.116 12.8525 ;
 RECT 73.892 12.6525 73.948 12.8525 ;
 RECT 73.052 12.6525 73.108 12.8525 ;
 RECT 72.884 12.6525 72.94 12.8525 ;
 RECT 73.388 12.6525 73.444 12.8525 ;
 RECT 73.22 12.6525 73.276 12.8525 ;
 RECT 72.38 12.6525 72.436 12.8525 ;
 RECT 72.212 12.6525 72.268 12.8525 ;
 RECT 72.716 12.6525 72.772 12.8525 ;
 RECT 72.548 12.6525 72.604 12.8525 ;
 RECT 71.708 12.6525 71.764 12.8525 ;
 RECT 71.54 12.6525 71.596 12.8525 ;
 RECT 72.044 12.6525 72.1 12.8525 ;
 RECT 71.876 12.6525 71.932 12.8525 ;
 RECT 71.036 12.6525 71.092 12.8525 ;
 RECT 70.868 12.6525 70.924 12.8525 ;
 RECT 71.372 12.6525 71.428 12.8525 ;
 RECT 71.204 12.6525 71.26 12.8525 ;
 RECT 70.364 12.6525 70.42 12.8525 ;
 RECT 70.7 12.6525 70.756 12.8525 ;
 RECT 70.532 12.6525 70.588 12.8525 ;
 RECT 74.732 14.4275 74.788 14.6275 ;
 RECT 74.06 14.4275 74.116 14.6275 ;
 RECT 73.388 14.4275 73.444 14.6275 ;
 RECT 72.716 14.4275 72.772 14.6275 ;
 RECT 72.044 14.4275 72.1 14.6275 ;
 RECT 71.372 14.4275 71.428 14.6275 ;
 RECT 70.7 14.4275 70.756 14.6275 ;
 END
 END vss.gds1225
 PIN vss.gds1226
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 17.782 0.29 17.982 ;
 END
 END vss.gds1226
 PIN vss.gds1227
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 19.057 2.962 19.257 ;
 END
 END vss.gds1227
 PIN vss.gds1228
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 20.317 2.962 20.517 ;
 END
 END vss.gds1228
 PIN vss.gds1229
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 19.482 0.602 19.682 ;
 END
 END vss.gds1229
 PIN vss.gds1230
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 17.683 0.942 17.883 ;
 END
 END vss.gds1230
 PIN vss.gds1231
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.646 16.884 1.702 17.084 ;
 END
 END vss.gds1231
 PIN vss.gds1232
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 19.065 1.282 19.265 ;
 END
 END vss.gds1232
 PIN vss.gds1233
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 17.987 2.122 18.187 ;
 END
 END vss.gds1233
 PIN vss.gds1234
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.754 17.4275 3.794 17.6275 ;
 END
 END vss.gds1234
 PIN vss.gds1235
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 17.5825 5.074 17.7825 ;
 END
 END vss.gds1235
 PIN vss.gds1236
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.282 16.274 4.338 16.474 ;
 END
 END vss.gds1236
 PIN vss.gds1237
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 18.1745 4.194 18.3745 ;
 END
 END vss.gds1237
 PIN vss.gds1238
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 19.916 3.142 20.116 ;
 END
 END vss.gds1238
 PIN vss.gds1239
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 20.099 4.882 20.299 ;
 END
 END vss.gds1239
 PIN vss.gds1240
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 17.607 4.002 17.807 ;
 END
 END vss.gds1240
 PIN vss.gds1241
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 17.7835 5.282 17.9835 ;
 END
 END vss.gds1241
 PIN vss.gds1242
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 17.516 2.302 17.716 ;
 END
 END vss.gds1242
 PIN vss.gds1243
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 16.739 3.142 16.939 ;
 END
 END vss.gds1243
 PIN vss.gds1244
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 19.202 1.462 19.402 ;
 END
 END vss.gds1244
 PIN vss.gds1245
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 17.76 0.718 17.96 ;
 END
 END vss.gds1245
 PIN vss.gds1246
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 3.5 18.512 3.556 18.663 ;
 RECT 3.248 18.491 3.304 18.663 ;
 RECT 4.004 18.512 4.06 18.663 ;
 RECT 3.752 18.491 3.808 18.663 ;
 RECT 1.568 17.386 1.624 17.586 ;
 RECT 0.98 17.386 1.036 17.586 ;
 RECT 2.996 17.386 3.052 17.586 ;
 RECT 3.248 17.246 3.304 17.446 ;
 RECT 3.5 17.2445 3.556 17.4445 ;
 RECT 4.088 17.246 4.144 17.446 ;
 RECT 3.92 17.246 3.976 17.446 ;
 RECT 1.988 17.106 2.044 17.306 ;
 RECT 2.996 17.106 3.052 17.306 ;
 RECT 3.5 16.023 3.556 16.205 ;
 RECT 0.56 16.023 0.616 16.223 ;
 RECT 1.568 16.023 1.624 16.223 ;
 RECT 0.98 16.023 1.036 16.223 ;
 RECT 2.576 16.023 2.632 16.223 ;
 RECT 2.156 16.023 2.212 16.223 ;
 RECT 1.988 16.023 2.044 16.223 ;
 RECT 3.248 15.902 3.304 16.102 ;
 RECT 3.5 15.799 3.556 15.981 ;
 RECT 4.088 15.902 4.144 16.102 ;
 RECT 3.92 15.902 3.976 16.102 ;
 RECT 2.576 19.0575 2.632 19.2575 ;
 RECT 2.408 19.0575 2.464 19.2575 ;
 RECT 2.996 19.0575 3.052 19.2575 ;
 RECT 3.332 19.149 3.388 19.349 ;
 RECT 3.5 19.1055 3.556 19.3055 ;
 RECT 0.98 18.9725 1.036 19.1725 ;
 RECT 2.072 18.973 2.128 19.173 ;
 RECT 2.576 20.3175 2.632 20.5175 ;
 RECT 2.408 20.3175 2.464 20.5175 ;
 RECT 2.996 20.3175 3.052 20.5175 ;
 RECT 3.332 20.409 3.388 20.609 ;
 RECT 3.5 20.3655 3.556 20.5655 ;
 RECT 0.98 20.2325 1.036 20.4325 ;
 RECT 2.072 20.233 2.128 20.433 ;
 RECT 0.392 20.323 0.448 20.523 ;
 RECT 0.812 20.409 0.868 20.609 ;
 RECT 0.644 20.323 0.7 20.523 ;
 RECT 1.232 20.323 1.288 20.523 ;
 RECT 1.4 20.323 1.456 20.523 ;
 RECT 1.568 20.323 1.624 20.523 ;
 RECT 1.82 20.323 1.876 20.523 ;
 RECT 2.24 20.323 2.296 20.523 ;
 RECT 2.744 20.233 2.8 20.433 ;
 RECT 3.164 20.323 3.22 20.523 ;
 RECT 3.92 20.323 3.976 20.523 ;
 RECT 0.392 19.063 0.448 19.263 ;
 RECT 0.812 19.149 0.868 19.349 ;
 RECT 0.644 19.063 0.7 19.263 ;
 RECT 1.232 19.063 1.288 19.263 ;
 RECT 1.4 19.063 1.456 19.263 ;
 RECT 1.568 19.063 1.624 19.263 ;
 RECT 1.82 19.063 1.876 19.263 ;
 RECT 2.24 19.063 2.296 19.263 ;
 RECT 2.744 18.973 2.8 19.173 ;
 RECT 3.164 19.063 3.22 19.263 ;
 RECT 3.92 19.063 3.976 19.263 ;
 RECT 3.752 19.333 3.808 19.533 ;
 RECT 4.508 19.2625 4.564 19.4625 ;
 RECT 2.156 17.125 2.212 17.325 ;
 RECT 0.56 17.086 0.616 17.286 ;
 RECT 1.568 17.0355 1.624 17.2355 ;
 RECT 0.98 17.0355 1.036 17.2355 ;
 RECT 0.56 15.6915 0.616 15.8915 ;
 RECT 1.568 15.6915 1.624 15.8915 ;
 RECT 0.98 15.6915 1.036 15.8915 ;
 RECT 2.072 15.762 2.128 15.962 ;
 RECT 1.904 15.762 1.96 15.962 ;
 RECT 3.08 15.762 3.136 15.962 ;
 RECT 2.912 15.762 2.968 15.962 ;
 RECT 2.744 15.762 2.8 15.962 ;
 RECT 4.676 15.902 4.732 16.102 ;
 RECT 4.424 15.8965 4.48 16.0965 ;
 RECT 0.56 17.367 0.616 17.567 ;
 RECT 2.408 17.265 2.464 17.465 ;
 RECT 2.24 17.367 2.296 17.567 ;
 RECT 2.072 17.367 2.128 17.567 ;
 RECT 2.744 17.246 2.8 17.446 ;
 RECT 4.676 17.246 4.732 17.446 ;
 RECT 4.424 17.246 4.48 17.446 ;
 RECT 0.56 18.469 0.616 18.669 ;
 RECT 1.568 18.469 1.624 18.669 ;
 RECT 0.98 18.469 1.036 18.669 ;
 RECT 1.988 18.448 2.044 18.648 ;
 RECT 2.492 18.448 2.548 18.648 ;
 RECT 2.24 18.448 2.296 18.648 ;
 RECT 2.744 18.448 2.8 18.648 ;
 RECT 2.996 18.448 3.052 18.648 ;
 RECT 4.676 18.448 4.732 18.648 ;
 RECT 4.424 18.448 4.48 18.648 ;
 END
 END vss.gds1246
 PIN vss.gds1247
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.046 15.902 10.086 16.102 ;
 END
 END vss.gds1247
 PIN vss.gds1248
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.374 15.902 9.414 16.102 ;
 END
 END vss.gds1248
 PIN vss.gds1249
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.702 15.902 8.742 16.102 ;
 END
 END vss.gds1249
 PIN vss.gds1250
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.03 15.902 8.07 16.102 ;
 END
 END vss.gds1250
 PIN vss.gds1251
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.778 15.695 9.824 15.895 ;
 END
 END vss.gds1251
 PIN vss.gds1252
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.174 15.695 10.214 15.895 ;
 END
 END vss.gds1252
 PIN vss.gds1253
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.106 15.695 9.152 15.895 ;
 END
 END vss.gds1253
 PIN vss.gds1254
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.502 15.695 9.542 15.895 ;
 END
 END vss.gds1254
 PIN vss.gds1255
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.434 15.695 8.48 15.895 ;
 END
 END vss.gds1255
 PIN vss.gds1256
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.83 15.695 8.87 15.895 ;
 END
 END vss.gds1256
 PIN vss.gds1257
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.762 15.695 7.808 15.895 ;
 END
 END vss.gds1257
 PIN vss.gds1258
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.158 15.695 8.198 15.895 ;
 END
 END vss.gds1258
 PIN vss.gds1259
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 18.1735 9.69 18.3735 ;
 END
 END vss.gds1259
 PIN vss.gds1260
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 18.1735 8.346 18.3735 ;
 END
 END vss.gds1260
 PIN vss.gds1261
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 18.1735 9.018 18.3735 ;
 END
 END vss.gds1261
 PIN vss.gds1262
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.942 16.8335 7.002 17.0335 ;
 END
 END vss.gds1262
 PIN vss.gds1263
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.09 15.695 7.136 15.895 ;
 END
 END vss.gds1263
 PIN vss.gds1264
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 18.1735 7.674 18.3735 ;
 END
 END vss.gds1264
 PIN vss.gds1265
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.358 15.902 7.398 16.102 ;
 END
 END vss.gds1265
 PIN vss.gds1266
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.486 15.695 7.526 15.895 ;
 END
 END vss.gds1266
 PIN vss.gds1267
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 17.5825 5.474 17.7825 ;
 END
 END vss.gds1267
 PIN vss.gds1268
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 17.5825 5.986 17.7825 ;
 END
 END vss.gds1268
 PIN vss.gds1269
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.734 16.9105 6.774 17.1105 ;
 END
 END vss.gds1269
 PIN vss.gds1270
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.606 16.9105 6.646 17.1105 ;
 END
 END vss.gds1270
 PIN vss.gds1271
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 17.999 6.178 18.199 ;
 END
 END vss.gds1271
 PIN vss.gds1272
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 17.6785 5.73 17.8785 ;
 END
 END vss.gds1272
 PIN vss.gds1273
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 18.246 6.434 18.446 ;
 END
 END vss.gds1273
 PIN vss.gds1274
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 10.136 18.493 10.192 18.693 ;
 RECT 9.632 18.483 9.688 18.683 ;
 RECT 9.464 18.493 9.52 18.693 ;
 RECT 8.96 18.483 9.016 18.683 ;
 RECT 8.792 18.493 8.848 18.693 ;
 RECT 8.288 18.483 8.344 18.683 ;
 RECT 8.12 18.493 8.176 18.693 ;
 RECT 6.944 18.483 7 18.683 ;
 RECT 7.616 18.483 7.672 18.683 ;
 RECT 7.448 18.493 7.504 18.693 ;
 RECT 5.6 17.386 5.656 17.586 ;
 RECT 9.968 15.721 10.024 15.921 ;
 RECT 9.8 15.721 9.856 15.921 ;
 RECT 10.136 15.736 10.192 15.936 ;
 RECT 9.296 15.721 9.352 15.921 ;
 RECT 9.128 15.721 9.184 15.921 ;
 RECT 9.464 15.736 9.52 15.936 ;
 RECT 9.632 15.736 9.688 15.936 ;
 RECT 8.624 15.721 8.68 15.921 ;
 RECT 8.456 15.721 8.512 15.921 ;
 RECT 8.792 15.736 8.848 15.936 ;
 RECT 8.96 15.736 9.016 15.936 ;
 RECT 7.952 15.721 8.008 15.921 ;
 RECT 7.784 15.721 7.84 15.921 ;
 RECT 8.12 15.736 8.176 15.936 ;
 RECT 8.288 15.736 8.344 15.936 ;
 RECT 7.28 15.721 7.336 15.921 ;
 RECT 7.112 15.721 7.168 15.921 ;
 RECT 6.944 15.736 7 15.936 ;
 RECT 7.448 15.736 7.504 15.936 ;
 RECT 7.616 15.736 7.672 15.936 ;
 RECT 9.968 16.795 10.024 16.995 ;
 RECT 9.8 16.795 9.856 16.995 ;
 RECT 10.136 16.795 10.192 16.995 ;
 RECT 9.296 16.795 9.352 16.995 ;
 RECT 9.128 16.795 9.184 16.995 ;
 RECT 9.632 16.795 9.688 16.995 ;
 RECT 9.464 16.795 9.52 16.995 ;
 RECT 8.624 16.795 8.68 16.995 ;
 RECT 8.456 16.795 8.512 16.995 ;
 RECT 8.96 16.795 9.016 16.995 ;
 RECT 8.792 16.795 8.848 16.995 ;
 RECT 7.952 16.795 8.008 16.995 ;
 RECT 7.784 16.795 7.84 16.995 ;
 RECT 8.288 16.795 8.344 16.995 ;
 RECT 8.12 16.795 8.176 16.995 ;
 RECT 7.28 16.795 7.336 16.995 ;
 RECT 6.944 16.795 7 16.995 ;
 RECT 7.112 16.795 7.168 16.995 ;
 RECT 7.616 16.795 7.672 16.995 ;
 RECT 7.448 16.795 7.504 16.995 ;
 RECT 6.524 20.285 6.58 20.485 ;
 RECT 6.524 19.025 6.58 19.225 ;
 RECT 6.692 19.348 6.748 19.548 ;
 RECT 6.608 19.333 6.664 19.533 ;
 RECT 5.432 15.902 5.488 16.102 ;
 RECT 5.6 15.902 5.656 16.102 ;
 RECT 5.768 15.902 5.824 16.102 ;
 RECT 5.936 15.902 5.992 16.102 ;
 RECT 6.44 15.902 6.496 16.102 ;
 RECT 6.104 15.902 6.16 16.102 ;
 RECT 6.272 15.902 6.328 16.102 ;
 RECT 5.432 17.246 5.488 17.446 ;
 RECT 5.6 17.106 5.656 17.306 ;
 RECT 5.768 17.246 5.824 17.446 ;
 RECT 5.936 17.246 5.992 17.446 ;
 RECT 6.104 17.246 6.16 17.446 ;
 RECT 6.272 17.246 6.328 17.446 ;
 RECT 6.44 17.246 6.496 17.446 ;
 RECT 5.432 18.448 5.488 18.648 ;
 RECT 5.6 18.448 5.656 18.648 ;
 RECT 5.768 18.448 5.824 18.648 ;
 RECT 5.936 18.448 5.992 18.648 ;
 RECT 6.104 18.448 6.16 18.648 ;
 RECT 6.272 18.448 6.328 18.648 ;
 RECT 6.44 18.448 6.496 18.648 ;
 END
 END vss.gds1274
 PIN vss.gds1275
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 19.602 14.87 19.802 ;
 END
 END vss.gds1275
 PIN vss.gds1276
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.262 16.9105 14.318 17.1105 ;
 END
 END vss.gds1276
 PIN vss.gds1277
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.062 15.902 12.102 16.102 ;
 END
 END vss.gds1277
 PIN vss.gds1278
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.39 15.902 11.43 16.102 ;
 END
 END vss.gds1278
 PIN vss.gds1279
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.718 15.902 10.758 16.102 ;
 END
 END vss.gds1279
 PIN vss.gds1280
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.794 15.695 11.84 15.895 ;
 END
 END vss.gds1280
 PIN vss.gds1281
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.19 15.695 12.23 15.895 ;
 END
 END vss.gds1281
 PIN vss.gds1282
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.122 15.695 11.168 15.895 ;
 END
 END vss.gds1282
 PIN vss.gds1283
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.518 15.695 11.558 15.895 ;
 END
 END vss.gds1283
 PIN vss.gds1284
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.45 15.695 10.496 15.895 ;
 END
 END vss.gds1284
 PIN vss.gds1285
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.846 15.695 10.886 15.895 ;
 END
 END vss.gds1285
 PIN vss.gds1286
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 16.3795 13.898 16.5795 ;
 END
 END vss.gds1286
 PIN vss.gds1287
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 16.1965 14.87 16.3965 ;
 END
 END vss.gds1287
 PIN vss.gds1288
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 18.2085 13.658 18.4085 ;
 END
 END vss.gds1288
 PIN vss.gds1289
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 16.022 13.058 16.222 ;
 END
 END vss.gds1289
 PIN vss.gds1290
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.262 19.151 13.318 19.351 ;
 END
 END vss.gds1290
 PIN vss.gds1291
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 18.1735 11.706 18.3735 ;
 END
 END vss.gds1291
 PIN vss.gds1292
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 18.1735 11.034 18.3735 ;
 END
 END vss.gds1292
 PIN vss.gds1293
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 18.3615 15.162 18.5615 ;
 END
 END vss.gds1293
 PIN vss.gds1294
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 18.1735 10.362 18.3735 ;
 END
 END vss.gds1294
 PIN vss.gds1295
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 18.4225 14.498 18.6225 ;
 END
 END vss.gds1295
 PIN vss.gds1296
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 18.3175 12.818 18.5175 ;
 END
 END vss.gds1296
 PIN vss.gds1297
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 17.757 12.378 17.957 ;
 END
 END vss.gds1297
 PIN vss.gds1298
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 17.5825 12.59 17.7825 ;
 END
 END vss.gds1298
 PIN vss.gds1299
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 19.562 13.898 19.762 ;
 END
 END vss.gds1299
 PIN vss.gds1300
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 13.244 18.389 13.3 18.589 ;
 RECT 12.32 18.483 12.376 18.683 ;
 RECT 12.152 18.493 12.208 18.693 ;
 RECT 11.648 18.483 11.704 18.683 ;
 RECT 11.48 18.493 11.536 18.693 ;
 RECT 10.976 18.483 11.032 18.683 ;
 RECT 10.808 18.493 10.864 18.693 ;
 RECT 10.304 18.483 10.36 18.683 ;
 RECT 12.824 16.042 12.88 16.242 ;
 RECT 15.176 16.042 15.232 16.242 ;
 RECT 15.008 16.042 15.064 16.242 ;
 RECT 13.664 16.023 13.72 16.223 ;
 RECT 12.992 16.023 13.048 16.223 ;
 RECT 13.16 16.023 13.216 16.223 ;
 RECT 13.496 16.023 13.552 16.223 ;
 RECT 14 16.023 14.056 16.223 ;
 RECT 14.168 16.023 14.224 16.223 ;
 RECT 13.832 16.023 13.888 16.223 ;
 RECT 14.84 16.023 14.896 16.223 ;
 RECT 14.504 16.042 14.56 16.242 ;
 RECT 14.672 16.042 14.728 16.242 ;
 RECT 13.244 15.762 13.3 15.962 ;
 RECT 13.58 15.762 13.636 15.962 ;
 RECT 12.908 15.762 12.964 15.962 ;
 RECT 13.916 15.762 13.972 15.962 ;
 RECT 14.252 15.762 14.308 15.962 ;
 RECT 14.924 15.762 14.98 15.962 ;
 RECT 11.984 15.721 12.04 15.921 ;
 RECT 11.816 15.721 11.872 15.921 ;
 RECT 12.152 15.736 12.208 15.936 ;
 RECT 12.32 15.736 12.376 15.936 ;
 RECT 11.312 15.721 11.368 15.921 ;
 RECT 11.144 15.721 11.2 15.921 ;
 RECT 11.48 15.736 11.536 15.936 ;
 RECT 11.648 15.736 11.704 15.936 ;
 RECT 10.64 15.721 10.696 15.921 ;
 RECT 10.472 15.721 10.528 15.921 ;
 RECT 10.808 15.736 10.864 15.936 ;
 RECT 10.976 15.736 11.032 15.936 ;
 RECT 10.304 15.736 10.36 15.936 ;
 RECT 14 19.74 14.056 19.913 ;
 RECT 14.168 19.713 14.224 19.913 ;
 RECT 14.336 20.333 14.392 20.533 ;
 RECT 14.168 20.333 14.224 20.533 ;
 RECT 13.16 17.379 13.216 17.579 ;
 RECT 13.412 17.593 13.468 17.793 ;
 RECT 11.984 16.795 12.04 16.995 ;
 RECT 11.816 16.795 11.872 16.995 ;
 RECT 12.32 16.795 12.376 16.995 ;
 RECT 12.152 16.795 12.208 16.995 ;
 RECT 11.312 16.795 11.368 16.995 ;
 RECT 11.144 16.795 11.2 16.995 ;
 RECT 11.648 16.795 11.704 16.995 ;
 RECT 11.48 16.795 11.536 16.995 ;
 RECT 10.64 16.795 10.696 16.995 ;
 RECT 10.472 16.795 10.528 16.995 ;
 RECT 10.976 16.795 11.032 16.995 ;
 RECT 10.808 16.795 10.864 16.995 ;
 RECT 10.304 16.795 10.36 16.995 ;
 RECT 14.336 19.073 14.392 19.273 ;
 RECT 14.168 19.073 14.224 19.273 ;
 RECT 15.008 19.283 15.064 19.483 ;
 RECT 14.84 19.757 14.896 19.922 ;
 RECT 14.672 19.757 14.728 19.922 ;
 RECT 13.664 19.207 13.72 19.407 ;
 END
 END vss.gds1300
 PIN vss.gds1301
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 20.317 16.146 20.517 ;
 END
 END vss.gds1301
 PIN vss.gds1302
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.958 15.902 19.998 16.102 ;
 END
 END vss.gds1302
 PIN vss.gds1303
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.286 15.902 19.326 16.102 ;
 END
 END vss.gds1303
 PIN vss.gds1304
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.614 15.902 18.654 16.102 ;
 END
 END vss.gds1304
 PIN vss.gds1305
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.69 15.695 19.736 15.895 ;
 END
 END vss.gds1305
 PIN vss.gds1306
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.086 15.695 20.126 15.895 ;
 END
 END vss.gds1306
 PIN vss.gds1307
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.018 15.695 19.064 15.895 ;
 END
 END vss.gds1307
 PIN vss.gds1308
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.414 15.695 19.454 15.895 ;
 END
 END vss.gds1308
 PIN vss.gds1309
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.346 15.695 18.392 15.895 ;
 END
 END vss.gds1309
 PIN vss.gds1310
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.742 15.695 18.782 15.895 ;
 END
 END vss.gds1310
 PIN vss.gds1311
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 16.1965 16.146 16.3965 ;
 END
 END vss.gds1311
 PIN vss.gds1312
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 20.117 15.418 20.317 ;
 END
 END vss.gds1312
 PIN vss.gds1313
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.438 18.943 17.494 19.143 ;
 END
 END vss.gds1313
 PIN vss.gds1314
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 18.1735 20.274 18.3735 ;
 END
 END vss.gds1314
 PIN vss.gds1315
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 16.44 16.814 16.64 ;
 END
 END vss.gds1315
 PIN vss.gds1316
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 19.9885 17.314 20.1885 ;
 END
 END vss.gds1316
 PIN vss.gds1317
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 18.1735 19.602 18.3735 ;
 END
 END vss.gds1317
 PIN vss.gds1318
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 18.1735 18.93 18.3735 ;
 END
 END vss.gds1318
 PIN vss.gds1319
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 18.144 16.994 18.344 ;
 END
 END vss.gds1319
 PIN vss.gds1320
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 18.4225 15.842 18.6225 ;
 END
 END vss.gds1320
 PIN vss.gds1321
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 18.3175 17.834 18.5175 ;
 END
 END vss.gds1321
 PIN vss.gds1322
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 18.197 16.49 18.397 ;
 END
 END vss.gds1322
 PIN vss.gds1323
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 19.057 16.146 19.257 ;
 END
 END vss.gds1323
 PIN vss.gds1324
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 17.757 18.258 17.957 ;
 END
 END vss.gds1324
 PIN vss.gds1325
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 20.216 18.483 20.272 18.683 ;
 RECT 20.048 18.493 20.104 18.693 ;
 RECT 19.544 18.483 19.6 18.683 ;
 RECT 19.376 18.493 19.432 18.693 ;
 RECT 18.2 18.483 18.256 18.683 ;
 RECT 18.872 18.483 18.928 18.683 ;
 RECT 18.704 18.493 18.76 18.693 ;
 RECT 16.1 16.042 16.156 16.242 ;
 RECT 15.596 16.042 15.652 16.242 ;
 RECT 15.428 16.042 15.484 16.242 ;
 RECT 15.764 16.042 15.82 16.242 ;
 RECT 16.604 16.042 16.66 16.242 ;
 RECT 16.772 16.042 16.828 16.242 ;
 RECT 16.436 16.042 16.492 16.242 ;
 RECT 16.268 16.042 16.324 16.242 ;
 RECT 17.696 16.042 17.752 16.242 ;
 RECT 17.276 16.023 17.332 16.205 ;
 RECT 17.024 16.023 17.08 16.205 ;
 RECT 19.88 15.721 19.936 15.921 ;
 RECT 19.712 15.721 19.768 15.921 ;
 RECT 20.048 15.736 20.104 15.936 ;
 RECT 20.216 15.736 20.272 15.936 ;
 RECT 15.26 15.762 15.316 15.962 ;
 RECT 15.596 15.762 15.652 15.962 ;
 RECT 15.932 15.762 15.988 15.962 ;
 RECT 16.268 15.762 16.324 15.962 ;
 RECT 17.192 15.799 17.248 15.981 ;
 RECT 16.94 15.799 16.996 15.981 ;
 RECT 17.528 15.762 17.584 15.962 ;
 RECT 17.78 15.762 17.836 15.962 ;
 RECT 19.208 15.721 19.264 15.921 ;
 RECT 19.04 15.721 19.096 15.921 ;
 RECT 19.376 15.736 19.432 15.936 ;
 RECT 19.544 15.736 19.6 15.936 ;
 RECT 18.2 15.736 18.256 15.936 ;
 RECT 18.704 15.736 18.76 15.936 ;
 RECT 18.872 15.736 18.928 15.936 ;
 RECT 15.596 18.724 15.652 18.924 ;
 RECT 15.848 18.727 15.904 18.927 ;
 RECT 16.52 19.76 16.576 19.913 ;
 RECT 15.764 19.757 15.82 19.922 ;
 RECT 15.596 19.757 15.652 19.922 ;
 RECT 15.596 19.984 15.652 20.184 ;
 RECT 15.848 19.987 15.904 20.187 ;
 RECT 18.536 15.721 18.592 15.921 ;
 RECT 18.368 15.721 18.424 15.921 ;
 RECT 18.116 16.574 18.172 16.774 ;
 RECT 19.88 16.795 19.936 16.995 ;
 RECT 19.712 16.795 19.768 16.995 ;
 RECT 20.216 16.795 20.272 16.995 ;
 RECT 20.048 16.795 20.104 16.995 ;
 RECT 19.208 16.795 19.264 16.995 ;
 RECT 19.04 16.795 19.096 16.995 ;
 RECT 19.544 16.795 19.6 16.995 ;
 RECT 19.376 16.795 19.432 16.995 ;
 RECT 18.536 16.795 18.592 16.995 ;
 RECT 18.2 16.795 18.256 16.995 ;
 RECT 18.368 16.795 18.424 16.995 ;
 RECT 18.872 16.795 18.928 16.995 ;
 RECT 18.704 16.795 18.76 16.995 ;
 RECT 16.856 20.3915 16.912 20.5915 ;
 RECT 15.428 19.283 15.484 19.483 ;
 RECT 16.352 19.3835 16.408 19.5835 ;
 RECT 16.856 19.1315 16.912 19.3315 ;
 END
 END vss.gds1325
 PIN vss.gds1326
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.082 15.902 25.122 16.102 ;
 END
 END vss.gds1326
 PIN vss.gds1327
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.41 15.902 24.45 16.102 ;
 END
 END vss.gds1327
 PIN vss.gds1328
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.318 15.902 23.358 16.102 ;
 END
 END vss.gds1328
 PIN vss.gds1329
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.646 15.902 22.686 16.102 ;
 END
 END vss.gds1329
 PIN vss.gds1330
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.974 15.902 22.014 16.102 ;
 END
 END vss.gds1330
 PIN vss.gds1331
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.302 15.902 21.342 16.102 ;
 END
 END vss.gds1331
 PIN vss.gds1332
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.63 15.902 20.67 16.102 ;
 END
 END vss.gds1332
 PIN vss.gds1333
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.814 15.695 24.86 15.895 ;
 END
 END vss.gds1333
 PIN vss.gds1334
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.21 15.695 25.25 15.895 ;
 END
 END vss.gds1334
 PIN vss.gds1335
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.142 15.695 24.188 15.895 ;
 END
 END vss.gds1335
 PIN vss.gds1336
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.538 15.695 24.578 15.895 ;
 END
 END vss.gds1336
 PIN vss.gds1337
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.05 15.695 23.096 15.895 ;
 END
 END vss.gds1337
 PIN vss.gds1338
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.446 15.695 23.486 15.895 ;
 END
 END vss.gds1338
 PIN vss.gds1339
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.378 15.695 22.424 15.895 ;
 END
 END vss.gds1339
 PIN vss.gds1340
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.774 15.695 22.814 15.895 ;
 END
 END vss.gds1340
 PIN vss.gds1341
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.706 15.695 21.752 15.895 ;
 END
 END vss.gds1341
 PIN vss.gds1342
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.102 15.695 22.142 15.895 ;
 END
 END vss.gds1342
 PIN vss.gds1343
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.034 15.695 21.08 15.895 ;
 END
 END vss.gds1343
 PIN vss.gds1344
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.43 15.695 21.47 15.895 ;
 END
 END vss.gds1344
 PIN vss.gds1345
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.362 15.695 20.408 15.895 ;
 END
 END vss.gds1345
 PIN vss.gds1346
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.758 15.695 20.798 15.895 ;
 END
 END vss.gds1346
 PIN vss.gds1347
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 18.1735 24.726 18.3735 ;
 END
 END vss.gds1347
 PIN vss.gds1348
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 18.1735 22.962 18.3735 ;
 END
 END vss.gds1348
 PIN vss.gds1349
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 18.1735 22.29 18.3735 ;
 END
 END vss.gds1349
 PIN vss.gds1350
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 18.1735 21.618 18.3735 ;
 END
 END vss.gds1350
 PIN vss.gds1351
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 18.1735 20.946 18.3735 ;
 END
 END vss.gds1351
 PIN vss.gds1352
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.994 16.8335 24.054 17.0335 ;
 END
 END vss.gds1352
 PIN vss.gds1353
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.722 16.9105 23.762 17.1105 ;
 END
 END vss.gds1353
 PIN vss.gds1354
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.866 16.9105 23.906 17.1105 ;
 END
 END vss.gds1354
 PIN vss.gds1355
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 18.1735 23.634 18.3735 ;
 END
 END vss.gds1355
 PIN vss.gds1356
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 25.172 18.493 25.228 18.693 ;
 RECT 23.996 18.483 24.052 18.683 ;
 RECT 24.668 18.483 24.724 18.683 ;
 RECT 24.5 18.493 24.556 18.693 ;
 RECT 23.576 18.483 23.632 18.683 ;
 RECT 23.408 18.493 23.464 18.693 ;
 RECT 22.904 18.483 22.96 18.683 ;
 RECT 22.736 18.493 22.792 18.693 ;
 RECT 22.232 18.483 22.288 18.683 ;
 RECT 22.064 18.493 22.12 18.693 ;
 RECT 21.56 18.483 21.616 18.683 ;
 RECT 21.392 18.493 21.448 18.693 ;
 RECT 20.888 18.483 20.944 18.683 ;
 RECT 20.72 18.493 20.776 18.693 ;
 RECT 25.004 15.721 25.06 15.921 ;
 RECT 24.836 15.721 24.892 15.921 ;
 RECT 25.172 15.736 25.228 15.936 ;
 RECT 23.996 15.736 24.052 15.936 ;
 RECT 24.5 15.736 24.556 15.936 ;
 RECT 24.668 15.736 24.724 15.936 ;
 RECT 23.408 15.736 23.464 15.936 ;
 RECT 23.576 15.736 23.632 15.936 ;
 RECT 22.568 15.721 22.624 15.921 ;
 RECT 22.4 15.721 22.456 15.921 ;
 RECT 22.736 15.736 22.792 15.936 ;
 RECT 22.904 15.736 22.96 15.936 ;
 RECT 21.896 15.721 21.952 15.921 ;
 RECT 21.728 15.721 21.784 15.921 ;
 RECT 22.064 15.736 22.12 15.936 ;
 RECT 22.232 15.736 22.288 15.936 ;
 RECT 21.224 15.721 21.28 15.921 ;
 RECT 21.056 15.721 21.112 15.921 ;
 RECT 21.392 15.736 21.448 15.936 ;
 RECT 21.56 15.736 21.616 15.936 ;
 RECT 20.72 15.736 20.776 15.936 ;
 RECT 20.888 15.736 20.944 15.936 ;
 RECT 20.552 15.721 20.608 15.921 ;
 RECT 20.384 15.721 20.44 15.921 ;
 RECT 24.332 15.721 24.388 15.921 ;
 RECT 24.164 15.721 24.22 15.921 ;
 RECT 23.24 15.721 23.296 15.921 ;
 RECT 23.072 15.721 23.128 15.921 ;
 RECT 25.004 16.795 25.06 16.995 ;
 RECT 24.836 16.795 24.892 16.995 ;
 RECT 25.172 16.795 25.228 16.995 ;
 RECT 24.332 16.795 24.388 16.995 ;
 RECT 23.996 16.795 24.052 16.995 ;
 RECT 24.164 16.795 24.22 16.995 ;
 RECT 24.668 16.795 24.724 16.995 ;
 RECT 24.5 16.795 24.556 16.995 ;
 RECT 23.24 16.795 23.296 16.995 ;
 RECT 23.072 16.795 23.128 16.995 ;
 RECT 23.576 16.795 23.632 16.995 ;
 RECT 23.408 16.795 23.464 16.995 ;
 RECT 22.568 16.795 22.624 16.995 ;
 RECT 22.4 16.795 22.456 16.995 ;
 RECT 22.904 16.795 22.96 16.995 ;
 RECT 22.736 16.795 22.792 16.995 ;
 RECT 21.896 16.795 21.952 16.995 ;
 RECT 21.728 16.795 21.784 16.995 ;
 RECT 22.232 16.795 22.288 16.995 ;
 RECT 22.064 16.795 22.12 16.995 ;
 RECT 21.224 16.795 21.28 16.995 ;
 RECT 21.056 16.795 21.112 16.995 ;
 RECT 21.56 16.795 21.616 16.995 ;
 RECT 21.392 16.795 21.448 16.995 ;
 RECT 20.552 16.795 20.608 16.995 ;
 RECT 20.888 16.795 20.944 16.995 ;
 RECT 20.72 16.795 20.776 16.995 ;
 RECT 20.384 16.795 20.44 16.995 ;
 RECT 23.912 19.22 23.968 19.42 ;
 RECT 23.744 18.6485 23.8 18.8485 ;
 END
 END vss.gds1356
 PIN vss.gds1357
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.114 15.902 29.154 16.102 ;
 END
 END vss.gds1357
 PIN vss.gds1358
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.442 15.902 28.482 16.102 ;
 END
 END vss.gds1358
 PIN vss.gds1359
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.77 15.902 27.81 16.102 ;
 END
 END vss.gds1359
 PIN vss.gds1360
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.098 15.902 27.138 16.102 ;
 END
 END vss.gds1360
 PIN vss.gds1361
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.426 15.902 26.466 16.102 ;
 END
 END vss.gds1361
 PIN vss.gds1362
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.754 15.902 25.794 16.102 ;
 END
 END vss.gds1362
 PIN vss.gds1363
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.846 15.695 28.892 15.895 ;
 END
 END vss.gds1363
 PIN vss.gds1364
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.242 15.695 29.282 15.895 ;
 END
 END vss.gds1364
 PIN vss.gds1365
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.174 15.695 28.22 15.895 ;
 END
 END vss.gds1365
 PIN vss.gds1366
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.57 15.695 28.61 15.895 ;
 END
 END vss.gds1366
 PIN vss.gds1367
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.502 15.695 27.548 15.895 ;
 END
 END vss.gds1367
 PIN vss.gds1368
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.898 15.695 27.938 15.895 ;
 END
 END vss.gds1368
 PIN vss.gds1369
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.83 15.695 26.876 15.895 ;
 END
 END vss.gds1369
 PIN vss.gds1370
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.226 15.695 27.266 15.895 ;
 END
 END vss.gds1370
 PIN vss.gds1371
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.158 15.695 26.204 15.895 ;
 END
 END vss.gds1371
 PIN vss.gds1372
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.554 15.695 26.594 15.895 ;
 END
 END vss.gds1372
 PIN vss.gds1373
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.486 15.695 25.532 15.895 ;
 END
 END vss.gds1373
 PIN vss.gds1374
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.882 15.695 25.922 15.895 ;
 END
 END vss.gds1374
 PIN vss.gds1375
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 17.757 29.43 17.957 ;
 END
 END vss.gds1375
 PIN vss.gds1376
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 18.1735 28.758 18.3735 ;
 END
 END vss.gds1376
 PIN vss.gds1377
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 18.1735 28.086 18.3735 ;
 END
 END vss.gds1377
 PIN vss.gds1378
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 18.1735 27.414 18.3735 ;
 END
 END vss.gds1378
 PIN vss.gds1379
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 18.1735 26.742 18.3735 ;
 END
 END vss.gds1379
 PIN vss.gds1380
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 18.1735 26.07 18.3735 ;
 END
 END vss.gds1380
 PIN vss.gds1381
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 18.1735 25.398 18.3735 ;
 END
 END vss.gds1381
 PIN vss.gds1382
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 16.022 30.11 16.222 ;
 END
 END vss.gds1382
 PIN vss.gds1383
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 18.3175 29.87 18.5175 ;
 END
 END vss.gds1383
 PIN vss.gds1384
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 17.5825 29.642 17.7825 ;
 END
 END vss.gds1384
 PIN vss.gds1385
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.372 18.483 29.428 18.683 ;
 RECT 29.204 18.493 29.26 18.693 ;
 RECT 28.7 18.483 28.756 18.683 ;
 RECT 28.532 18.493 28.588 18.693 ;
 RECT 28.028 18.483 28.084 18.683 ;
 RECT 27.86 18.493 27.916 18.693 ;
 RECT 27.356 18.483 27.412 18.683 ;
 RECT 27.188 18.493 27.244 18.693 ;
 RECT 26.684 18.483 26.74 18.683 ;
 RECT 26.516 18.493 26.572 18.693 ;
 RECT 26.012 18.483 26.068 18.683 ;
 RECT 25.844 18.493 25.9 18.693 ;
 RECT 25.34 18.483 25.396 18.683 ;
 RECT 29.876 16.042 29.932 16.242 ;
 RECT 30.044 16.023 30.1 16.223 ;
 RECT 30.212 16.023 30.268 16.223 ;
 RECT 29.96 15.762 30.016 15.962 ;
 RECT 29.036 15.721 29.092 15.921 ;
 RECT 28.868 15.721 28.924 15.921 ;
 RECT 29.204 15.736 29.26 15.936 ;
 RECT 29.372 15.736 29.428 15.936 ;
 RECT 28.364 15.721 28.42 15.921 ;
 RECT 28.196 15.721 28.252 15.921 ;
 RECT 28.532 15.736 28.588 15.936 ;
 RECT 28.7 15.736 28.756 15.936 ;
 RECT 27.692 15.721 27.748 15.921 ;
 RECT 27.524 15.721 27.58 15.921 ;
 RECT 27.86 15.736 27.916 15.936 ;
 RECT 28.028 15.736 28.084 15.936 ;
 RECT 27.02 15.721 27.076 15.921 ;
 RECT 26.852 15.721 26.908 15.921 ;
 RECT 27.188 15.736 27.244 15.936 ;
 RECT 27.356 15.736 27.412 15.936 ;
 RECT 26.348 15.721 26.404 15.921 ;
 RECT 26.18 15.721 26.236 15.921 ;
 RECT 26.516 15.736 26.572 15.936 ;
 RECT 26.684 15.736 26.74 15.936 ;
 RECT 25.676 15.721 25.732 15.921 ;
 RECT 25.508 15.721 25.564 15.921 ;
 RECT 25.844 15.736 25.9 15.936 ;
 RECT 26.012 15.736 26.068 15.936 ;
 RECT 25.34 15.736 25.396 15.936 ;
 RECT 30.212 17.379 30.268 17.579 ;
 RECT 29.036 16.795 29.092 16.995 ;
 RECT 28.868 16.795 28.924 16.995 ;
 RECT 29.372 16.795 29.428 16.995 ;
 RECT 29.204 16.795 29.26 16.995 ;
 RECT 28.364 16.795 28.42 16.995 ;
 RECT 28.196 16.795 28.252 16.995 ;
 RECT 28.7 16.795 28.756 16.995 ;
 RECT 28.532 16.795 28.588 16.995 ;
 RECT 27.692 16.795 27.748 16.995 ;
 RECT 27.524 16.795 27.58 16.995 ;
 RECT 28.028 16.795 28.084 16.995 ;
 RECT 27.86 16.795 27.916 16.995 ;
 RECT 27.02 16.795 27.076 16.995 ;
 RECT 26.852 16.795 26.908 16.995 ;
 RECT 27.356 16.795 27.412 16.995 ;
 RECT 27.188 16.795 27.244 16.995 ;
 RECT 26.348 16.795 26.404 16.995 ;
 RECT 26.18 16.795 26.236 16.995 ;
 RECT 26.684 16.795 26.74 16.995 ;
 RECT 26.516 16.795 26.572 16.995 ;
 RECT 25.676 16.795 25.732 16.995 ;
 RECT 25.508 16.795 25.564 16.995 ;
 RECT 26.012 16.795 26.068 16.995 ;
 RECT 25.844 16.795 25.9 16.995 ;
 RECT 25.34 16.795 25.396 16.995 ;
 END
 END vss.gds1385
 PIN vss.gds1386
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 19.602 31.922 19.802 ;
 END
 END vss.gds1386
 PIN vss.gds1387
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 19.562 30.95 19.762 ;
 END
 END vss.gds1387
 PIN vss.gds1388
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.314 16.9105 31.37 17.1105 ;
 END
 END vss.gds1388
 PIN vss.gds1389
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 20.317 33.198 20.517 ;
 END
 END vss.gds1389
 PIN vss.gds1390
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 20.117 32.47 20.317 ;
 END
 END vss.gds1390
 PIN vss.gds1391
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 16.1965 31.922 16.3965 ;
 END
 END vss.gds1391
 PIN vss.gds1392
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 16.1965 33.198 16.3965 ;
 END
 END vss.gds1392
 PIN vss.gds1393
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.314 19.151 30.37 19.351 ;
 END
 END vss.gds1393
 PIN vss.gds1394
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 18.4225 32.894 18.6225 ;
 END
 END vss.gds1394
 PIN vss.gds1395
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 18.3615 32.214 18.5615 ;
 END
 END vss.gds1395
 PIN vss.gds1396
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.49 18.943 34.546 19.143 ;
 END
 END vss.gds1396
 PIN vss.gds1397
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 18.2085 30.71 18.4085 ;
 END
 END vss.gds1397
 PIN vss.gds1398
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 16.44 33.866 16.64 ;
 END
 END vss.gds1398
 PIN vss.gds1399
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 19.057 33.198 19.257 ;
 END
 END vss.gds1399
 PIN vss.gds1400
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 18.197 33.542 18.397 ;
 END
 END vss.gds1400
 PIN vss.gds1401
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 19.9885 34.366 20.1885 ;
 END
 END vss.gds1401
 PIN vss.gds1402
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 18.4225 31.55 18.6225 ;
 END
 END vss.gds1402
 PIN vss.gds1403
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 18.3175 34.886 18.5175 ;
 END
 END vss.gds1403
 PIN vss.gds1404
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 18.144 34.046 18.344 ;
 END
 END vss.gds1404
 PIN vss.gds1405
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 16.3795 30.95 16.5795 ;
 END
 END vss.gds1405
 PIN vss.gds1406
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 30.296 18.389 30.352 18.589 ;
 RECT 32.228 16.042 32.284 16.242 ;
 RECT 32.06 16.042 32.116 16.242 ;
 RECT 30.716 16.023 30.772 16.223 ;
 RECT 30.548 16.023 30.604 16.223 ;
 RECT 31.052 16.023 31.108 16.223 ;
 RECT 31.22 16.023 31.276 16.223 ;
 RECT 30.884 16.023 30.94 16.223 ;
 RECT 31.892 16.023 31.948 16.223 ;
 RECT 31.556 16.042 31.612 16.242 ;
 RECT 31.724 16.042 31.78 16.242 ;
 RECT 33.152 16.042 33.208 16.242 ;
 RECT 32.648 16.042 32.704 16.242 ;
 RECT 32.48 16.042 32.536 16.242 ;
 RECT 32.816 16.042 32.872 16.242 ;
 RECT 33.656 16.042 33.712 16.242 ;
 RECT 33.824 16.042 33.88 16.242 ;
 RECT 33.488 16.042 33.544 16.242 ;
 RECT 33.32 16.042 33.376 16.242 ;
 RECT 34.748 16.042 34.804 16.242 ;
 RECT 34.328 16.023 34.384 16.205 ;
 RECT 34.076 16.023 34.132 16.205 ;
 RECT 32.312 15.762 32.368 15.962 ;
 RECT 30.296 15.762 30.352 15.962 ;
 RECT 30.632 15.762 30.688 15.962 ;
 RECT 30.968 15.762 31.024 15.962 ;
 RECT 31.304 15.762 31.36 15.962 ;
 RECT 31.976 15.762 32.032 15.962 ;
 RECT 32.648 15.762 32.704 15.962 ;
 RECT 32.984 15.762 33.04 15.962 ;
 RECT 33.32 15.762 33.376 15.962 ;
 RECT 34.244 15.799 34.3 15.981 ;
 RECT 33.992 15.799 34.048 15.981 ;
 RECT 34.58 15.762 34.636 15.962 ;
 RECT 34.832 15.762 34.888 15.962 ;
 RECT 32.648 18.724 32.704 18.924 ;
 RECT 32.9 18.727 32.956 18.927 ;
 RECT 33.572 19.76 33.628 19.913 ;
 RECT 31.052 19.74 31.108 19.913 ;
 RECT 31.22 19.713 31.276 19.913 ;
 RECT 32.816 19.757 32.872 19.922 ;
 RECT 32.648 19.757 32.704 19.922 ;
 RECT 31.892 19.757 31.948 19.922 ;
 RECT 31.724 19.757 31.78 19.922 ;
 RECT 31.388 19.073 31.444 19.273 ;
 RECT 31.22 19.073 31.276 19.273 ;
 RECT 30.716 19.207 30.772 19.407 ;
 RECT 32.648 19.984 32.704 20.184 ;
 RECT 32.9 19.987 32.956 20.187 ;
 RECT 35.168 16.574 35.224 16.774 ;
 RECT 32.06 19.283 32.116 19.483 ;
 RECT 32.48 19.283 32.536 19.483 ;
 RECT 31.388 20.333 31.444 20.533 ;
 RECT 31.22 20.333 31.276 20.533 ;
 RECT 30.464 17.593 30.52 17.793 ;
 RECT 33.908 20.3915 33.964 20.5915 ;
 RECT 33.908 19.1315 33.964 19.3315 ;
 RECT 33.404 19.3835 33.46 19.5835 ;
 END
 END vss.gds1406
 PIN vss.gds1407
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.698 15.902 39.738 16.102 ;
 END
 END vss.gds1407
 PIN vss.gds1408
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.026 15.902 39.066 16.102 ;
 END
 END vss.gds1408
 PIN vss.gds1409
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.354 15.902 38.394 16.102 ;
 END
 END vss.gds1409
 PIN vss.gds1410
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.682 15.902 37.722 16.102 ;
 END
 END vss.gds1410
 PIN vss.gds1411
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.01 15.902 37.05 16.102 ;
 END
 END vss.gds1411
 PIN vss.gds1412
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.338 15.902 36.378 16.102 ;
 END
 END vss.gds1412
 PIN vss.gds1413
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.666 15.902 35.706 16.102 ;
 END
 END vss.gds1413
 PIN vss.gds1414
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.102 15.695 40.148 15.895 ;
 END
 END vss.gds1414
 PIN vss.gds1415
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.43 15.695 39.476 15.895 ;
 END
 END vss.gds1415
 PIN vss.gds1416
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.826 15.695 39.866 15.895 ;
 END
 END vss.gds1416
 PIN vss.gds1417
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.758 15.695 38.804 15.895 ;
 END
 END vss.gds1417
 PIN vss.gds1418
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.154 15.695 39.194 15.895 ;
 END
 END vss.gds1418
 PIN vss.gds1419
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.086 15.695 38.132 15.895 ;
 END
 END vss.gds1419
 PIN vss.gds1420
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.482 15.695 38.522 15.895 ;
 END
 END vss.gds1420
 PIN vss.gds1421
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.414 15.695 37.46 15.895 ;
 END
 END vss.gds1421
 PIN vss.gds1422
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.81 15.695 37.85 15.895 ;
 END
 END vss.gds1422
 PIN vss.gds1423
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.742 15.695 36.788 15.895 ;
 END
 END vss.gds1423
 PIN vss.gds1424
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.138 15.695 37.178 15.895 ;
 END
 END vss.gds1424
 PIN vss.gds1425
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.07 15.695 36.116 15.895 ;
 END
 END vss.gds1425
 PIN vss.gds1426
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.466 15.695 36.506 15.895 ;
 END
 END vss.gds1426
 PIN vss.gds1427
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.398 15.695 35.444 15.895 ;
 END
 END vss.gds1427
 PIN vss.gds1428
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.794 15.695 35.834 15.895 ;
 END
 END vss.gds1428
 PIN vss.gds1429
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 18.1735 37.998 18.3735 ;
 END
 END vss.gds1429
 PIN vss.gds1430
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 18.1735 37.326 18.3735 ;
 END
 END vss.gds1430
 PIN vss.gds1431
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 18.1735 38.67 18.3735 ;
 END
 END vss.gds1431
 PIN vss.gds1432
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 18.1735 36.654 18.3735 ;
 END
 END vss.gds1432
 PIN vss.gds1433
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 18.1735 39.342 18.3735 ;
 END
 END vss.gds1433
 PIN vss.gds1434
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 18.1735 40.014 18.3735 ;
 END
 END vss.gds1434
 PIN vss.gds1435
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 17.757 35.31 17.957 ;
 END
 END vss.gds1435
 PIN vss.gds1436
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 18.1735 35.982 18.3735 ;
 END
 END vss.gds1436
 PIN vss.gds1437
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 39.956 18.483 40.012 18.683 ;
 RECT 39.788 18.493 39.844 18.693 ;
 RECT 39.284 18.483 39.34 18.683 ;
 RECT 39.116 18.493 39.172 18.693 ;
 RECT 38.612 18.483 38.668 18.683 ;
 RECT 38.444 18.493 38.5 18.693 ;
 RECT 37.94 18.483 37.996 18.683 ;
 RECT 37.772 18.493 37.828 18.693 ;
 RECT 37.268 18.483 37.324 18.683 ;
 RECT 37.1 18.493 37.156 18.693 ;
 RECT 36.596 18.483 36.652 18.683 ;
 RECT 36.428 18.493 36.484 18.693 ;
 RECT 35.252 18.483 35.308 18.683 ;
 RECT 35.924 18.483 35.98 18.683 ;
 RECT 35.756 18.493 35.812 18.693 ;
 RECT 39.62 15.721 39.676 15.921 ;
 RECT 39.452 15.721 39.508 15.921 ;
 RECT 39.788 15.736 39.844 15.936 ;
 RECT 39.956 15.736 40.012 15.936 ;
 RECT 38.948 15.721 39.004 15.921 ;
 RECT 38.78 15.721 38.836 15.921 ;
 RECT 39.116 15.736 39.172 15.936 ;
 RECT 39.284 15.736 39.34 15.936 ;
 RECT 38.276 15.721 38.332 15.921 ;
 RECT 38.108 15.721 38.164 15.921 ;
 RECT 38.444 15.736 38.5 15.936 ;
 RECT 38.612 15.736 38.668 15.936 ;
 RECT 37.604 15.721 37.66 15.921 ;
 RECT 37.436 15.721 37.492 15.921 ;
 RECT 37.772 15.736 37.828 15.936 ;
 RECT 37.94 15.736 37.996 15.936 ;
 RECT 36.932 15.721 36.988 15.921 ;
 RECT 36.764 15.721 36.82 15.921 ;
 RECT 37.1 15.736 37.156 15.936 ;
 RECT 37.268 15.736 37.324 15.936 ;
 RECT 36.26 15.721 36.316 15.921 ;
 RECT 36.092 15.721 36.148 15.921 ;
 RECT 36.428 15.736 36.484 15.936 ;
 RECT 36.596 15.736 36.652 15.936 ;
 RECT 35.252 15.736 35.308 15.936 ;
 RECT 35.756 15.736 35.812 15.936 ;
 RECT 35.924 15.736 35.98 15.936 ;
 RECT 40.124 15.721 40.18 15.921 ;
 RECT 35.588 15.721 35.644 15.921 ;
 RECT 35.42 15.721 35.476 15.921 ;
 RECT 40.124 16.795 40.18 16.995 ;
 RECT 39.62 16.795 39.676 16.995 ;
 RECT 39.452 16.795 39.508 16.995 ;
 RECT 39.956 16.795 40.012 16.995 ;
 RECT 39.788 16.795 39.844 16.995 ;
 RECT 38.948 16.795 39.004 16.995 ;
 RECT 38.78 16.795 38.836 16.995 ;
 RECT 39.284 16.795 39.34 16.995 ;
 RECT 39.116 16.795 39.172 16.995 ;
 RECT 38.276 16.795 38.332 16.995 ;
 RECT 38.108 16.795 38.164 16.995 ;
 RECT 38.612 16.795 38.668 16.995 ;
 RECT 38.444 16.795 38.5 16.995 ;
 RECT 37.604 16.795 37.66 16.995 ;
 RECT 37.436 16.795 37.492 16.995 ;
 RECT 37.94 16.795 37.996 16.995 ;
 RECT 37.772 16.795 37.828 16.995 ;
 RECT 36.932 16.795 36.988 16.995 ;
 RECT 36.764 16.795 36.82 16.995 ;
 RECT 37.268 16.795 37.324 16.995 ;
 RECT 37.1 16.795 37.156 16.995 ;
 RECT 36.26 16.795 36.316 16.995 ;
 RECT 36.092 16.795 36.148 16.995 ;
 RECT 36.596 16.795 36.652 16.995 ;
 RECT 36.428 16.795 36.484 16.995 ;
 RECT 35.588 16.795 35.644 16.995 ;
 RECT 35.252 16.795 35.308 16.995 ;
 RECT 35.42 16.795 35.476 16.995 ;
 RECT 35.924 16.795 35.98 16.995 ;
 RECT 35.756 16.795 35.812 16.995 ;
 END
 END vss.gds1437
 PIN vss.gds1438
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.822 15.902 44.862 16.102 ;
 END
 END vss.gds1438
 PIN vss.gds1439
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.15 15.902 44.19 16.102 ;
 END
 END vss.gds1439
 PIN vss.gds1440
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.478 15.902 43.518 16.102 ;
 END
 END vss.gds1440
 PIN vss.gds1441
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.806 15.902 42.846 16.102 ;
 END
 END vss.gds1441
 PIN vss.gds1442
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.134 15.902 42.174 16.102 ;
 END
 END vss.gds1442
 PIN vss.gds1443
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.462 15.902 41.502 16.102 ;
 END
 END vss.gds1443
 PIN vss.gds1444
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.37 15.902 40.41 16.102 ;
 END
 END vss.gds1444
 PIN vss.gds1445
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.226 15.695 45.272 15.895 ;
 END
 END vss.gds1445
 PIN vss.gds1446
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.554 15.695 44.6 15.895 ;
 END
 END vss.gds1446
 PIN vss.gds1447
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.95 15.695 44.99 15.895 ;
 END
 END vss.gds1447
 PIN vss.gds1448
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.882 15.695 43.928 15.895 ;
 END
 END vss.gds1448
 PIN vss.gds1449
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.278 15.695 44.318 15.895 ;
 END
 END vss.gds1449
 PIN vss.gds1450
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.21 15.695 43.256 15.895 ;
 END
 END vss.gds1450
 PIN vss.gds1451
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.606 15.695 43.646 15.895 ;
 END
 END vss.gds1451
 PIN vss.gds1452
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.538 15.695 42.584 15.895 ;
 END
 END vss.gds1452
 PIN vss.gds1453
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.934 15.695 42.974 15.895 ;
 END
 END vss.gds1453
 PIN vss.gds1454
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.866 15.695 41.912 15.895 ;
 END
 END vss.gds1454
 PIN vss.gds1455
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.262 15.695 42.302 15.895 ;
 END
 END vss.gds1455
 PIN vss.gds1456
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.194 15.695 41.24 15.895 ;
 END
 END vss.gds1456
 PIN vss.gds1457
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.59 15.695 41.63 15.895 ;
 END
 END vss.gds1457
 PIN vss.gds1458
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.498 15.695 40.538 15.895 ;
 END
 END vss.gds1458
 PIN vss.gds1459
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.774 16.9105 40.814 17.1105 ;
 END
 END vss.gds1459
 PIN vss.gds1460
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.918 16.9105 40.958 17.1105 ;
 END
 END vss.gds1460
 PIN vss.gds1461
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 18.1735 45.138 18.3735 ;
 END
 END vss.gds1461
 PIN vss.gds1462
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 18.1735 44.466 18.3735 ;
 END
 END vss.gds1462
 PIN vss.gds1463
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 18.1735 43.794 18.3735 ;
 END
 END vss.gds1463
 PIN vss.gds1464
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 18.1735 43.122 18.3735 ;
 END
 END vss.gds1464
 PIN vss.gds1465
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 18.1735 42.45 18.3735 ;
 END
 END vss.gds1465
 PIN vss.gds1466
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 18.1735 41.778 18.3735 ;
 END
 END vss.gds1466
 PIN vss.gds1467
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 18.1735 40.686 18.3735 ;
 END
 END vss.gds1467
 PIN vss.gds1468
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.046 16.8335 41.106 17.0335 ;
 END
 END vss.gds1468
 PIN vss.gds1469
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 45.08 18.483 45.136 18.683 ;
 RECT 44.912 18.493 44.968 18.693 ;
 RECT 44.408 18.483 44.464 18.683 ;
 RECT 44.24 18.493 44.296 18.693 ;
 RECT 43.736 18.483 43.792 18.683 ;
 RECT 43.568 18.493 43.624 18.693 ;
 RECT 43.064 18.483 43.12 18.683 ;
 RECT 42.896 18.493 42.952 18.693 ;
 RECT 42.392 18.483 42.448 18.683 ;
 RECT 42.224 18.493 42.28 18.693 ;
 RECT 41.048 18.483 41.104 18.683 ;
 RECT 41.72 18.483 41.776 18.683 ;
 RECT 41.552 18.493 41.608 18.693 ;
 RECT 40.628 18.483 40.684 18.683 ;
 RECT 40.46 18.493 40.516 18.693 ;
 RECT 44.744 15.721 44.8 15.921 ;
 RECT 44.576 15.721 44.632 15.921 ;
 RECT 44.912 15.736 44.968 15.936 ;
 RECT 45.08 15.736 45.136 15.936 ;
 RECT 44.072 15.721 44.128 15.921 ;
 RECT 43.904 15.721 43.96 15.921 ;
 RECT 44.24 15.736 44.296 15.936 ;
 RECT 44.408 15.736 44.464 15.936 ;
 RECT 43.4 15.721 43.456 15.921 ;
 RECT 43.232 15.721 43.288 15.921 ;
 RECT 43.568 15.736 43.624 15.936 ;
 RECT 43.736 15.736 43.792 15.936 ;
 RECT 42.728 15.721 42.784 15.921 ;
 RECT 42.56 15.721 42.616 15.921 ;
 RECT 42.896 15.736 42.952 15.936 ;
 RECT 43.064 15.736 43.12 15.936 ;
 RECT 42.056 15.721 42.112 15.921 ;
 RECT 41.888 15.721 41.944 15.921 ;
 RECT 42.224 15.736 42.28 15.936 ;
 RECT 42.392 15.736 42.448 15.936 ;
 RECT 41.048 15.736 41.104 15.936 ;
 RECT 41.552 15.736 41.608 15.936 ;
 RECT 41.72 15.736 41.776 15.936 ;
 RECT 40.46 15.736 40.516 15.936 ;
 RECT 40.628 15.736 40.684 15.936 ;
 RECT 41.384 15.721 41.44 15.921 ;
 RECT 41.216 15.721 41.272 15.921 ;
 RECT 40.292 15.721 40.348 15.921 ;
 RECT 44.744 16.795 44.8 16.995 ;
 RECT 44.576 16.795 44.632 16.995 ;
 RECT 45.08 16.795 45.136 16.995 ;
 RECT 44.912 16.795 44.968 16.995 ;
 RECT 44.072 16.795 44.128 16.995 ;
 RECT 43.904 16.795 43.96 16.995 ;
 RECT 44.408 16.795 44.464 16.995 ;
 RECT 44.24 16.795 44.296 16.995 ;
 RECT 43.4 16.795 43.456 16.995 ;
 RECT 43.232 16.795 43.288 16.995 ;
 RECT 43.736 16.795 43.792 16.995 ;
 RECT 43.568 16.795 43.624 16.995 ;
 RECT 42.728 16.795 42.784 16.995 ;
 RECT 42.56 16.795 42.616 16.995 ;
 RECT 43.064 16.795 43.12 16.995 ;
 RECT 42.896 16.795 42.952 16.995 ;
 RECT 42.056 16.795 42.112 16.995 ;
 RECT 41.888 16.795 41.944 16.995 ;
 RECT 42.392 16.795 42.448 16.995 ;
 RECT 42.224 16.795 42.28 16.995 ;
 RECT 41.384 16.795 41.44 16.995 ;
 RECT 41.048 16.795 41.104 16.995 ;
 RECT 41.216 16.795 41.272 16.995 ;
 RECT 41.72 16.795 41.776 16.995 ;
 RECT 41.552 16.795 41.608 16.995 ;
 RECT 40.628 16.795 40.684 16.995 ;
 RECT 40.46 16.795 40.516 16.995 ;
 RECT 40.292 16.795 40.348 16.995 ;
 RECT 40.964 19.22 41.02 19.42 ;
 RECT 40.796 18.6485 40.852 18.8485 ;
 END
 END vss.gds1469
 PIN vss.gds1470
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 19.602 48.974 19.802 ;
 END
 END vss.gds1470
 PIN vss.gds1471
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 19.562 48.002 19.762 ;
 END
 END vss.gds1471
 PIN vss.gds1472
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.366 16.9105 48.422 17.1105 ;
 END
 END vss.gds1472
 PIN vss.gds1473
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 20.317 50.25 20.517 ;
 END
 END vss.gds1473
 PIN vss.gds1474
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.166 15.902 46.206 16.102 ;
 END
 END vss.gds1474
 PIN vss.gds1475
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.494 15.902 45.534 16.102 ;
 END
 END vss.gds1475
 PIN vss.gds1476
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.898 15.695 45.944 15.895 ;
 END
 END vss.gds1476
 PIN vss.gds1477
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.294 15.695 46.334 15.895 ;
 END
 END vss.gds1477
 PIN vss.gds1478
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.622 15.695 45.662 15.895 ;
 END
 END vss.gds1478
 PIN vss.gds1479
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 16.1965 48.974 16.3965 ;
 END
 END vss.gds1479
 PIN vss.gds1480
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 16.1965 50.25 16.3965 ;
 END
 END vss.gds1480
 PIN vss.gds1481
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 20.117 49.522 20.317 ;
 END
 END vss.gds1481
 PIN vss.gds1482
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.366 19.151 47.422 19.351 ;
 END
 END vss.gds1482
 PIN vss.gds1483
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 18.1735 45.81 18.3735 ;
 END
 END vss.gds1483
 PIN vss.gds1484
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 17.757 46.482 17.957 ;
 END
 END vss.gds1484
 PIN vss.gds1485
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 16.022 47.162 16.222 ;
 END
 END vss.gds1485
 PIN vss.gds1486
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 18.3175 46.922 18.5175 ;
 END
 END vss.gds1486
 PIN vss.gds1487
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 16.3795 48.002 16.5795 ;
 END
 END vss.gds1487
 PIN vss.gds1488
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 17.5825 46.694 17.7825 ;
 END
 END vss.gds1488
 PIN vss.gds1489
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 18.2085 47.762 18.4085 ;
 END
 END vss.gds1489
 PIN vss.gds1490
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 18.3615 49.266 18.5615 ;
 END
 END vss.gds1490
 PIN vss.gds1491
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 18.4225 48.602 18.6225 ;
 END
 END vss.gds1491
 PIN vss.gds1492
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 18.4225 49.946 18.6225 ;
 END
 END vss.gds1492
 PIN vss.gds1493
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 19.057 50.25 19.257 ;
 END
 END vss.gds1493
 PIN vss.gds1494
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 47.348 18.389 47.404 18.589 ;
 RECT 46.424 18.483 46.48 18.683 ;
 RECT 46.256 18.493 46.312 18.693 ;
 RECT 45.752 18.483 45.808 18.683 ;
 RECT 45.584 18.493 45.64 18.693 ;
 RECT 46.928 16.042 46.984 16.242 ;
 RECT 49.28 16.042 49.336 16.242 ;
 RECT 49.112 16.042 49.168 16.242 ;
 RECT 47.768 16.023 47.824 16.223 ;
 RECT 47.096 16.023 47.152 16.223 ;
 RECT 47.264 16.023 47.32 16.223 ;
 RECT 47.6 16.023 47.656 16.223 ;
 RECT 48.104 16.023 48.16 16.223 ;
 RECT 48.272 16.023 48.328 16.223 ;
 RECT 47.936 16.023 47.992 16.223 ;
 RECT 48.944 16.023 49 16.223 ;
 RECT 48.608 16.042 48.664 16.242 ;
 RECT 48.776 16.042 48.832 16.242 ;
 RECT 50.204 16.042 50.26 16.242 ;
 RECT 49.7 16.042 49.756 16.242 ;
 RECT 49.532 16.042 49.588 16.242 ;
 RECT 49.868 16.042 49.924 16.242 ;
 RECT 49.364 15.762 49.42 15.962 ;
 RECT 47.348 15.762 47.404 15.962 ;
 RECT 47.684 15.762 47.74 15.962 ;
 RECT 47.012 15.762 47.068 15.962 ;
 RECT 48.02 15.762 48.076 15.962 ;
 RECT 48.356 15.762 48.412 15.962 ;
 RECT 49.028 15.762 49.084 15.962 ;
 RECT 49.7 15.762 49.756 15.962 ;
 RECT 50.036 15.762 50.092 15.962 ;
 RECT 46.088 15.721 46.144 15.921 ;
 RECT 45.92 15.721 45.976 15.921 ;
 RECT 46.256 15.736 46.312 15.936 ;
 RECT 46.424 15.736 46.48 15.936 ;
 RECT 45.416 15.721 45.472 15.921 ;
 RECT 45.248 15.721 45.304 15.921 ;
 RECT 45.584 15.736 45.64 15.936 ;
 RECT 45.752 15.736 45.808 15.936 ;
 RECT 49.7 18.724 49.756 18.924 ;
 RECT 49.952 18.727 50.008 18.927 ;
 RECT 48.104 19.74 48.16 19.913 ;
 RECT 48.272 19.713 48.328 19.913 ;
 RECT 49.868 19.757 49.924 19.922 ;
 RECT 49.7 19.757 49.756 19.922 ;
 RECT 48.944 19.757 49 19.922 ;
 RECT 48.776 19.757 48.832 19.922 ;
 RECT 49.7 19.984 49.756 20.184 ;
 RECT 49.952 19.987 50.008 20.187 ;
 RECT 48.44 19.073 48.496 19.273 ;
 RECT 48.272 19.073 48.328 19.273 ;
 RECT 47.768 19.207 47.824 19.407 ;
 RECT 47.264 17.379 47.32 17.579 ;
 RECT 47.516 17.593 47.572 17.793 ;
 RECT 49.112 19.283 49.168 19.483 ;
 RECT 49.532 19.283 49.588 19.483 ;
 RECT 48.44 20.333 48.496 20.533 ;
 RECT 48.272 20.333 48.328 20.533 ;
 RECT 46.088 16.795 46.144 16.995 ;
 RECT 45.92 16.795 45.976 16.995 ;
 RECT 46.424 16.795 46.48 16.995 ;
 RECT 46.256 16.795 46.312 16.995 ;
 RECT 45.416 16.795 45.472 16.995 ;
 RECT 45.248 16.795 45.304 16.995 ;
 RECT 45.752 16.795 45.808 16.995 ;
 RECT 45.584 16.795 45.64 16.995 ;
 END
 END vss.gds1494
 PIN vss.gds1495
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.734 15.902 54.774 16.102 ;
 END
 END vss.gds1495
 PIN vss.gds1496
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.062 15.902 54.102 16.102 ;
 END
 END vss.gds1496
 PIN vss.gds1497
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.39 15.902 53.43 16.102 ;
 END
 END vss.gds1497
 PIN vss.gds1498
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.718 15.902 52.758 16.102 ;
 END
 END vss.gds1498
 PIN vss.gds1499
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.138 15.695 55.184 15.895 ;
 END
 END vss.gds1499
 PIN vss.gds1500
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.466 15.695 54.512 15.895 ;
 END
 END vss.gds1500
 PIN vss.gds1501
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.862 15.695 54.902 15.895 ;
 END
 END vss.gds1501
 PIN vss.gds1502
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.794 15.695 53.84 15.895 ;
 END
 END vss.gds1502
 PIN vss.gds1503
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.19 15.695 54.23 15.895 ;
 END
 END vss.gds1503
 PIN vss.gds1504
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.122 15.695 53.168 15.895 ;
 END
 END vss.gds1504
 PIN vss.gds1505
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.518 15.695 53.558 15.895 ;
 END
 END vss.gds1505
 PIN vss.gds1506
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.45 15.695 52.496 15.895 ;
 END
 END vss.gds1506
 PIN vss.gds1507
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.846 15.695 52.886 15.895 ;
 END
 END vss.gds1507
 PIN vss.gds1508
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 18.1735 54.378 18.3735 ;
 END
 END vss.gds1508
 PIN vss.gds1509
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 18.1735 55.05 18.3735 ;
 END
 END vss.gds1509
 PIN vss.gds1510
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 16.44 50.918 16.64 ;
 END
 END vss.gds1510
 PIN vss.gds1511
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.542 18.943 51.598 19.143 ;
 END
 END vss.gds1511
 PIN vss.gds1512
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 18.1735 53.706 18.3735 ;
 END
 END vss.gds1512
 PIN vss.gds1513
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 19.9885 51.418 20.1885 ;
 END
 END vss.gds1513
 PIN vss.gds1514
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 18.1735 53.034 18.3735 ;
 END
 END vss.gds1514
 PIN vss.gds1515
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 18.3175 51.938 18.5175 ;
 END
 END vss.gds1515
 PIN vss.gds1516
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 18.197 50.594 18.397 ;
 END
 END vss.gds1516
 PIN vss.gds1517
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 17.757 52.362 17.957 ;
 END
 END vss.gds1517
 PIN vss.gds1518
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 18.144 51.098 18.344 ;
 END
 END vss.gds1518
 PIN vss.gds1519
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 54.992 18.483 55.048 18.683 ;
 RECT 54.824 18.493 54.88 18.693 ;
 RECT 54.32 18.483 54.376 18.683 ;
 RECT 54.152 18.493 54.208 18.693 ;
 RECT 53.648 18.483 53.704 18.683 ;
 RECT 53.48 18.493 53.536 18.693 ;
 RECT 52.304 18.483 52.36 18.683 ;
 RECT 52.976 18.483 53.032 18.683 ;
 RECT 52.808 18.493 52.864 18.693 ;
 RECT 50.708 16.042 50.764 16.242 ;
 RECT 50.876 16.042 50.932 16.242 ;
 RECT 50.54 16.042 50.596 16.242 ;
 RECT 50.372 16.042 50.428 16.242 ;
 RECT 51.8 16.042 51.856 16.242 ;
 RECT 51.38 16.023 51.436 16.205 ;
 RECT 51.128 16.023 51.184 16.205 ;
 RECT 55.16 15.721 55.216 15.921 ;
 RECT 54.656 15.721 54.712 15.921 ;
 RECT 54.488 15.721 54.544 15.921 ;
 RECT 54.824 15.736 54.88 15.936 ;
 RECT 54.992 15.736 55.048 15.936 ;
 RECT 53.984 15.721 54.04 15.921 ;
 RECT 53.816 15.721 53.872 15.921 ;
 RECT 54.152 15.736 54.208 15.936 ;
 RECT 54.32 15.736 54.376 15.936 ;
 RECT 50.372 15.762 50.428 15.962 ;
 RECT 51.296 15.799 51.352 15.981 ;
 RECT 51.044 15.799 51.1 15.981 ;
 RECT 51.632 15.762 51.688 15.962 ;
 RECT 51.884 15.762 51.94 15.962 ;
 RECT 53.312 15.721 53.368 15.921 ;
 RECT 53.144 15.721 53.2 15.921 ;
 RECT 53.48 15.736 53.536 15.936 ;
 RECT 53.648 15.736 53.704 15.936 ;
 RECT 52.304 15.736 52.36 15.936 ;
 RECT 52.808 15.736 52.864 15.936 ;
 RECT 52.976 15.736 53.032 15.936 ;
 RECT 50.624 19.76 50.68 19.913 ;
 RECT 52.22 16.574 52.276 16.774 ;
 RECT 52.64 15.721 52.696 15.921 ;
 RECT 52.472 15.721 52.528 15.921 ;
 RECT 55.16 16.795 55.216 16.995 ;
 RECT 54.656 16.795 54.712 16.995 ;
 RECT 54.488 16.795 54.544 16.995 ;
 RECT 54.992 16.795 55.048 16.995 ;
 RECT 54.824 16.795 54.88 16.995 ;
 RECT 53.984 16.795 54.04 16.995 ;
 RECT 53.816 16.795 53.872 16.995 ;
 RECT 54.32 16.795 54.376 16.995 ;
 RECT 54.152 16.795 54.208 16.995 ;
 RECT 53.312 16.795 53.368 16.995 ;
 RECT 53.144 16.795 53.2 16.995 ;
 RECT 53.648 16.795 53.704 16.995 ;
 RECT 53.48 16.795 53.536 16.995 ;
 RECT 52.64 16.795 52.696 16.995 ;
 RECT 52.304 16.795 52.36 16.995 ;
 RECT 52.472 16.795 52.528 16.995 ;
 RECT 52.976 16.795 53.032 16.995 ;
 RECT 52.808 16.795 52.864 16.995 ;
 RECT 50.96 20.3915 51.016 20.5915 ;
 RECT 50.456 19.3835 50.512 19.5835 ;
 RECT 50.96 19.1315 51.016 19.3315 ;
 END
 END vss.gds1519
 PIN vss.gds1520
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.858 15.902 59.898 16.102 ;
 END
 END vss.gds1520
 PIN vss.gds1521
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.186 15.902 59.226 16.102 ;
 END
 END vss.gds1521
 PIN vss.gds1522
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.514 15.902 58.554 16.102 ;
 END
 END vss.gds1522
 PIN vss.gds1523
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.422 15.902 57.462 16.102 ;
 END
 END vss.gds1523
 PIN vss.gds1524
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.75 15.902 56.79 16.102 ;
 END
 END vss.gds1524
 PIN vss.gds1525
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.078 15.902 56.118 16.102 ;
 END
 END vss.gds1525
 PIN vss.gds1526
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.406 15.902 55.446 16.102 ;
 END
 END vss.gds1526
 PIN vss.gds1527
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.59 15.695 59.636 15.895 ;
 END
 END vss.gds1527
 PIN vss.gds1528
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.986 15.695 60.026 15.895 ;
 END
 END vss.gds1528
 PIN vss.gds1529
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.918 15.695 58.964 15.895 ;
 END
 END vss.gds1529
 PIN vss.gds1530
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.314 15.695 59.354 15.895 ;
 END
 END vss.gds1530
 PIN vss.gds1531
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.246 15.695 58.292 15.895 ;
 END
 END vss.gds1531
 PIN vss.gds1532
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.642 15.695 58.682 15.895 ;
 END
 END vss.gds1532
 PIN vss.gds1533
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.154 15.695 57.2 15.895 ;
 END
 END vss.gds1533
 PIN vss.gds1534
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.55 15.695 57.59 15.895 ;
 END
 END vss.gds1534
 PIN vss.gds1535
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.482 15.695 56.528 15.895 ;
 END
 END vss.gds1535
 PIN vss.gds1536
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.878 15.695 56.918 15.895 ;
 END
 END vss.gds1536
 PIN vss.gds1537
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.81 15.695 55.856 15.895 ;
 END
 END vss.gds1537
 PIN vss.gds1538
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.206 15.695 56.246 15.895 ;
 END
 END vss.gds1538
 PIN vss.gds1539
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.534 15.695 55.574 15.895 ;
 END
 END vss.gds1539
 PIN vss.gds1540
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.826 16.9105 57.866 17.1105 ;
 END
 END vss.gds1540
 PIN vss.gds1541
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.97 16.9105 58.01 17.1105 ;
 END
 END vss.gds1541
 PIN vss.gds1542
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.098 16.8335 58.158 17.0335 ;
 END
 END vss.gds1542
 PIN vss.gds1543
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 18.1735 60.174 18.3735 ;
 END
 END vss.gds1543
 PIN vss.gds1544
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 18.1735 59.502 18.3735 ;
 END
 END vss.gds1544
 PIN vss.gds1545
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 18.1735 58.83 18.3735 ;
 END
 END vss.gds1545
 PIN vss.gds1546
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 18.1735 55.722 18.3735 ;
 END
 END vss.gds1546
 PIN vss.gds1547
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 18.1735 56.394 18.3735 ;
 END
 END vss.gds1547
 PIN vss.gds1548
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 18.1735 57.738 18.3735 ;
 END
 END vss.gds1548
 PIN vss.gds1549
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 18.1735 57.066 18.3735 ;
 END
 END vss.gds1549
 PIN vss.gds1550
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 60.116 18.483 60.172 18.683 ;
 RECT 59.948 18.493 60.004 18.693 ;
 RECT 59.444 18.483 59.5 18.683 ;
 RECT 59.276 18.493 59.332 18.693 ;
 RECT 58.1 18.483 58.156 18.683 ;
 RECT 58.772 18.483 58.828 18.683 ;
 RECT 58.604 18.493 58.66 18.693 ;
 RECT 57.68 18.483 57.736 18.683 ;
 RECT 57.512 18.493 57.568 18.693 ;
 RECT 57.008 18.483 57.064 18.683 ;
 RECT 56.84 18.493 56.896 18.693 ;
 RECT 56.336 18.483 56.392 18.683 ;
 RECT 56.168 18.493 56.224 18.693 ;
 RECT 55.664 18.483 55.72 18.683 ;
 RECT 55.496 18.493 55.552 18.693 ;
 RECT 59.78 15.721 59.836 15.921 ;
 RECT 59.612 15.721 59.668 15.921 ;
 RECT 59.948 15.736 60.004 15.936 ;
 RECT 60.116 15.736 60.172 15.936 ;
 RECT 59.108 15.721 59.164 15.921 ;
 RECT 58.94 15.721 58.996 15.921 ;
 RECT 59.276 15.736 59.332 15.936 ;
 RECT 59.444 15.736 59.5 15.936 ;
 RECT 58.1 15.736 58.156 15.936 ;
 RECT 58.604 15.736 58.66 15.936 ;
 RECT 58.772 15.736 58.828 15.936 ;
 RECT 57.512 15.736 57.568 15.936 ;
 RECT 57.68 15.736 57.736 15.936 ;
 RECT 56.672 15.721 56.728 15.921 ;
 RECT 56.504 15.721 56.56 15.921 ;
 RECT 56.84 15.736 56.896 15.936 ;
 RECT 57.008 15.736 57.064 15.936 ;
 RECT 56 15.721 56.056 15.921 ;
 RECT 55.832 15.721 55.888 15.921 ;
 RECT 56.168 15.736 56.224 15.936 ;
 RECT 56.336 15.736 56.392 15.936 ;
 RECT 55.328 15.721 55.384 15.921 ;
 RECT 55.496 15.736 55.552 15.936 ;
 RECT 55.664 15.736 55.72 15.936 ;
 RECT 58.436 15.721 58.492 15.921 ;
 RECT 58.268 15.721 58.324 15.921 ;
 RECT 57.344 15.721 57.4 15.921 ;
 RECT 57.176 15.721 57.232 15.921 ;
 RECT 59.78 16.795 59.836 16.995 ;
 RECT 59.612 16.795 59.668 16.995 ;
 RECT 60.116 16.795 60.172 16.995 ;
 RECT 59.948 16.795 60.004 16.995 ;
 RECT 59.108 16.795 59.164 16.995 ;
 RECT 58.94 16.795 58.996 16.995 ;
 RECT 59.444 16.795 59.5 16.995 ;
 RECT 59.276 16.795 59.332 16.995 ;
 RECT 58.436 16.795 58.492 16.995 ;
 RECT 58.1 16.795 58.156 16.995 ;
 RECT 58.268 16.795 58.324 16.995 ;
 RECT 58.772 16.795 58.828 16.995 ;
 RECT 58.604 16.795 58.66 16.995 ;
 RECT 57.344 16.795 57.4 16.995 ;
 RECT 57.176 16.795 57.232 16.995 ;
 RECT 57.68 16.795 57.736 16.995 ;
 RECT 57.512 16.795 57.568 16.995 ;
 RECT 56.672 16.795 56.728 16.995 ;
 RECT 56.504 16.795 56.56 16.995 ;
 RECT 57.008 16.795 57.064 16.995 ;
 RECT 56.84 16.795 56.896 16.995 ;
 RECT 56 16.795 56.056 16.995 ;
 RECT 55.832 16.795 55.888 16.995 ;
 RECT 56.336 16.795 56.392 16.995 ;
 RECT 56.168 16.795 56.224 16.995 ;
 RECT 55.328 16.795 55.384 16.995 ;
 RECT 55.664 16.795 55.72 16.995 ;
 RECT 55.496 16.795 55.552 16.995 ;
 RECT 58.016 19.22 58.072 19.42 ;
 RECT 57.848 18.6485 57.904 18.8485 ;
 END
 END vss.gds1550
 PIN vss.gds1551
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 19.562 65.054 19.762 ;
 END
 END vss.gds1551
 PIN vss.gds1552
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.218 15.902 63.258 16.102 ;
 END
 END vss.gds1552
 PIN vss.gds1553
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.546 15.902 62.586 16.102 ;
 END
 END vss.gds1553
 PIN vss.gds1554
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.874 15.902 61.914 16.102 ;
 END
 END vss.gds1554
 PIN vss.gds1555
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.202 15.902 61.242 16.102 ;
 END
 END vss.gds1555
 PIN vss.gds1556
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.53 15.902 60.57 16.102 ;
 END
 END vss.gds1556
 PIN vss.gds1557
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.95 15.695 62.996 15.895 ;
 END
 END vss.gds1557
 PIN vss.gds1558
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.346 15.695 63.386 15.895 ;
 END
 END vss.gds1558
 PIN vss.gds1559
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.278 15.695 62.324 15.895 ;
 END
 END vss.gds1559
 PIN vss.gds1560
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.674 15.695 62.714 15.895 ;
 END
 END vss.gds1560
 PIN vss.gds1561
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.606 15.695 61.652 15.895 ;
 END
 END vss.gds1561
 PIN vss.gds1562
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.002 15.695 62.042 15.895 ;
 END
 END vss.gds1562
 PIN vss.gds1563
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.934 15.695 60.98 15.895 ;
 END
 END vss.gds1563
 PIN vss.gds1564
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.33 15.695 61.37 15.895 ;
 END
 END vss.gds1564
 PIN vss.gds1565
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.262 15.695 60.308 15.895 ;
 END
 END vss.gds1565
 PIN vss.gds1566
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.658 15.695 60.698 15.895 ;
 END
 END vss.gds1566
 PIN vss.gds1567
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 16.022 64.214 16.222 ;
 END
 END vss.gds1567
 PIN vss.gds1568
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.418 19.151 64.474 19.351 ;
 END
 END vss.gds1568
 PIN vss.gds1569
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 17.757 63.534 17.957 ;
 END
 END vss.gds1569
 PIN vss.gds1570
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 18.1735 62.862 18.3735 ;
 END
 END vss.gds1570
 PIN vss.gds1571
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 18.1735 62.19 18.3735 ;
 END
 END vss.gds1571
 PIN vss.gds1572
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 18.1735 61.518 18.3735 ;
 END
 END vss.gds1572
 PIN vss.gds1573
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 18.1735 60.846 18.3735 ;
 END
 END vss.gds1573
 PIN vss.gds1574
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 18.3175 63.974 18.5175 ;
 END
 END vss.gds1574
 PIN vss.gds1575
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 16.3795 65.054 16.5795 ;
 END
 END vss.gds1575
 PIN vss.gds1576
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 17.5825 63.746 17.7825 ;
 END
 END vss.gds1576
 PIN vss.gds1577
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 18.2085 64.814 18.4085 ;
 END
 END vss.gds1577
 PIN vss.gds1578
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 64.4 18.389 64.456 18.589 ;
 RECT 63.476 18.483 63.532 18.683 ;
 RECT 63.308 18.493 63.364 18.693 ;
 RECT 62.804 18.483 62.86 18.683 ;
 RECT 62.636 18.493 62.692 18.693 ;
 RECT 62.132 18.483 62.188 18.683 ;
 RECT 61.964 18.493 62.02 18.693 ;
 RECT 61.46 18.483 61.516 18.683 ;
 RECT 61.292 18.493 61.348 18.693 ;
 RECT 60.788 18.483 60.844 18.683 ;
 RECT 60.62 18.493 60.676 18.693 ;
 RECT 63.98 16.042 64.036 16.242 ;
 RECT 64.82 16.023 64.876 16.223 ;
 RECT 64.148 16.023 64.204 16.223 ;
 RECT 64.316 16.023 64.372 16.223 ;
 RECT 64.652 16.023 64.708 16.223 ;
 RECT 65.156 16.023 65.212 16.223 ;
 RECT 64.988 16.023 65.044 16.223 ;
 RECT 64.4 15.762 64.456 15.962 ;
 RECT 64.736 15.762 64.792 15.962 ;
 RECT 64.064 15.762 64.12 15.962 ;
 RECT 65.072 15.762 65.128 15.962 ;
 RECT 63.14 15.721 63.196 15.921 ;
 RECT 62.972 15.721 63.028 15.921 ;
 RECT 63.308 15.736 63.364 15.936 ;
 RECT 63.476 15.736 63.532 15.936 ;
 RECT 62.468 15.721 62.524 15.921 ;
 RECT 62.3 15.721 62.356 15.921 ;
 RECT 62.636 15.736 62.692 15.936 ;
 RECT 62.804 15.736 62.86 15.936 ;
 RECT 61.796 15.721 61.852 15.921 ;
 RECT 61.628 15.721 61.684 15.921 ;
 RECT 61.964 15.736 62.02 15.936 ;
 RECT 62.132 15.736 62.188 15.936 ;
 RECT 61.124 15.721 61.18 15.921 ;
 RECT 60.956 15.721 61.012 15.921 ;
 RECT 61.292 15.736 61.348 15.936 ;
 RECT 61.46 15.736 61.516 15.936 ;
 RECT 60.62 15.736 60.676 15.936 ;
 RECT 60.788 15.736 60.844 15.936 ;
 RECT 60.452 15.721 60.508 15.921 ;
 RECT 60.284 15.721 60.34 15.921 ;
 RECT 65.156 19.74 65.212 19.913 ;
 RECT 64.82 19.207 64.876 19.407 ;
 RECT 64.316 17.379 64.372 17.579 ;
 RECT 64.568 17.593 64.624 17.793 ;
 RECT 63.14 16.795 63.196 16.995 ;
 RECT 62.972 16.795 63.028 16.995 ;
 RECT 63.476 16.795 63.532 16.995 ;
 RECT 63.308 16.795 63.364 16.995 ;
 RECT 62.468 16.795 62.524 16.995 ;
 RECT 62.3 16.795 62.356 16.995 ;
 RECT 62.804 16.795 62.86 16.995 ;
 RECT 62.636 16.795 62.692 16.995 ;
 RECT 61.796 16.795 61.852 16.995 ;
 RECT 61.628 16.795 61.684 16.995 ;
 RECT 62.132 16.795 62.188 16.995 ;
 RECT 61.964 16.795 62.02 16.995 ;
 RECT 61.124 16.795 61.18 16.995 ;
 RECT 60.956 16.795 61.012 16.995 ;
 RECT 61.46 16.795 61.516 16.995 ;
 RECT 61.292 16.795 61.348 16.995 ;
 RECT 60.452 16.795 60.508 16.995 ;
 RECT 60.788 16.795 60.844 16.995 ;
 RECT 60.62 16.795 60.676 16.995 ;
 RECT 60.284 16.795 60.34 16.995 ;
 END
 END vss.gds1578
 PIN vss.gds1579
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 19.602 66.026 19.802 ;
 END
 END vss.gds1579
 PIN vss.gds1580
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.418 16.9105 65.474 17.1105 ;
 END
 END vss.gds1580
 PIN vss.gds1581
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.77 15.902 69.81 16.102 ;
 END
 END vss.gds1581
 PIN vss.gds1582
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.174 15.695 70.22 15.895 ;
 END
 END vss.gds1582
 PIN vss.gds1583
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.502 15.695 69.548 15.895 ;
 END
 END vss.gds1583
 PIN vss.gds1584
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.898 15.695 69.938 15.895 ;
 END
 END vss.gds1584
 PIN vss.gds1585
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 16.1965 66.026 16.3965 ;
 END
 END vss.gds1585
 PIN vss.gds1586
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 16.1965 67.302 16.3965 ;
 END
 END vss.gds1586
 PIN vss.gds1587
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 20.317 67.302 20.517 ;
 END
 END vss.gds1587
 PIN vss.gds1588
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 18.3615 66.318 18.5615 ;
 END
 END vss.gds1588
 PIN vss.gds1589
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 20.117 66.574 20.317 ;
 END
 END vss.gds1589
 PIN vss.gds1590
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 18.1735 70.086 18.3735 ;
 END
 END vss.gds1590
 PIN vss.gds1591
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.594 18.943 68.65 19.143 ;
 END
 END vss.gds1591
 PIN vss.gds1592
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 16.44 67.97 16.64 ;
 END
 END vss.gds1592
 PIN vss.gds1593
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 18.144 68.15 18.344 ;
 END
 END vss.gds1593
 PIN vss.gds1594
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 19.9885 68.47 20.1885 ;
 END
 END vss.gds1594
 PIN vss.gds1595
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 19.057 67.302 19.257 ;
 END
 END vss.gds1595
 PIN vss.gds1596
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 18.197 67.646 18.397 ;
 END
 END vss.gds1596
 PIN vss.gds1597
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 18.4225 65.654 18.6225 ;
 END
 END vss.gds1597
 PIN vss.gds1598
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 18.4225 66.998 18.6225 ;
 END
 END vss.gds1598
 PIN vss.gds1599
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 18.3175 68.99 18.5175 ;
 END
 END vss.gds1599
 PIN vss.gds1600
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 17.757 69.414 17.957 ;
 END
 END vss.gds1600
 PIN vss.gds1601
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 69.356 18.483 69.412 18.683 ;
 RECT 70.028 18.483 70.084 18.683 ;
 RECT 69.86 18.493 69.916 18.693 ;
 RECT 66.332 16.042 66.388 16.242 ;
 RECT 66.164 16.042 66.22 16.242 ;
 RECT 65.324 16.023 65.38 16.223 ;
 RECT 65.996 16.023 66.052 16.223 ;
 RECT 65.66 16.042 65.716 16.242 ;
 RECT 65.828 16.042 65.884 16.242 ;
 RECT 67.256 16.042 67.312 16.242 ;
 RECT 66.752 16.042 66.808 16.242 ;
 RECT 66.584 16.042 66.64 16.242 ;
 RECT 66.92 16.042 66.976 16.242 ;
 RECT 67.76 16.042 67.816 16.242 ;
 RECT 67.928 16.042 67.984 16.242 ;
 RECT 67.592 16.042 67.648 16.242 ;
 RECT 67.424 16.042 67.48 16.242 ;
 RECT 68.852 16.042 68.908 16.242 ;
 RECT 68.432 16.023 68.488 16.205 ;
 RECT 68.18 16.023 68.236 16.205 ;
 RECT 66.416 15.762 66.472 15.962 ;
 RECT 65.408 15.762 65.464 15.962 ;
 RECT 66.08 15.762 66.136 15.962 ;
 RECT 66.752 15.762 66.808 15.962 ;
 RECT 67.088 15.762 67.144 15.962 ;
 RECT 67.424 15.762 67.48 15.962 ;
 RECT 68.348 15.799 68.404 15.981 ;
 RECT 68.096 15.799 68.152 15.981 ;
 RECT 68.684 15.762 68.74 15.962 ;
 RECT 68.936 15.762 68.992 15.962 ;
 RECT 70.196 15.721 70.252 15.921 ;
 RECT 69.356 15.736 69.412 15.936 ;
 RECT 69.86 15.736 69.916 15.936 ;
 RECT 70.028 15.736 70.084 15.936 ;
 RECT 66.752 18.724 66.808 18.924 ;
 RECT 67.004 18.727 67.06 18.927 ;
 RECT 67.676 19.76 67.732 19.913 ;
 RECT 65.324 19.713 65.38 19.913 ;
 RECT 66.92 19.757 66.976 19.922 ;
 RECT 66.752 19.757 66.808 19.922 ;
 RECT 65.996 19.757 66.052 19.922 ;
 RECT 65.828 19.757 65.884 19.922 ;
 RECT 66.752 19.984 66.808 20.184 ;
 RECT 67.004 19.987 67.06 20.187 ;
 RECT 65.492 19.073 65.548 19.273 ;
 RECT 65.324 19.073 65.38 19.273 ;
 RECT 69.692 15.721 69.748 15.921 ;
 RECT 69.524 15.721 69.58 15.921 ;
 RECT 69.272 16.574 69.328 16.774 ;
 RECT 66.164 19.283 66.22 19.483 ;
 RECT 66.584 19.283 66.64 19.483 ;
 RECT 65.492 20.333 65.548 20.533 ;
 RECT 65.324 20.333 65.38 20.533 ;
 RECT 68.012 20.3915 68.068 20.5915 ;
 RECT 67.508 19.3835 67.564 19.5835 ;
 RECT 68.012 19.1315 68.068 19.3315 ;
 RECT 70.196 16.795 70.252 16.995 ;
 RECT 69.692 16.795 69.748 16.995 ;
 RECT 69.356 16.795 69.412 16.995 ;
 RECT 69.524 16.795 69.58 16.995 ;
 RECT 70.028 16.795 70.084 16.995 ;
 RECT 69.86 16.795 69.916 16.995 ;
 END
 END vss.gds1601
 PIN vss.gds1602
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.474 15.902 74.514 16.102 ;
 END
 END vss.gds1602
 PIN vss.gds1603
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.802 15.902 73.842 16.102 ;
 END
 END vss.gds1603
 PIN vss.gds1604
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.13 15.902 73.17 16.102 ;
 END
 END vss.gds1604
 PIN vss.gds1605
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.458 15.902 72.498 16.102 ;
 END
 END vss.gds1605
 PIN vss.gds1606
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.786 15.902 71.826 16.102 ;
 END
 END vss.gds1606
 PIN vss.gds1607
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.114 15.902 71.154 16.102 ;
 END
 END vss.gds1607
 PIN vss.gds1608
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.442 15.902 70.482 16.102 ;
 END
 END vss.gds1608
 PIN vss.gds1609
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.206 15.695 74.252 15.895 ;
 END
 END vss.gds1609
 PIN vss.gds1610
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.602 15.695 74.642 15.895 ;
 END
 END vss.gds1610
 PIN vss.gds1611
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.534 15.695 73.58 15.895 ;
 END
 END vss.gds1611
 PIN vss.gds1612
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.93 15.695 73.97 15.895 ;
 END
 END vss.gds1612
 PIN vss.gds1613
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.862 15.695 72.908 15.895 ;
 END
 END vss.gds1613
 PIN vss.gds1614
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.258 15.695 73.298 15.895 ;
 END
 END vss.gds1614
 PIN vss.gds1615
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.19 15.695 72.236 15.895 ;
 END
 END vss.gds1615
 PIN vss.gds1616
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.586 15.695 72.626 15.895 ;
 END
 END vss.gds1616
 PIN vss.gds1617
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.518 15.695 71.564 15.895 ;
 END
 END vss.gds1617
 PIN vss.gds1618
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.914 15.695 71.954 15.895 ;
 END
 END vss.gds1618
 PIN vss.gds1619
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.846 15.695 70.892 15.895 ;
 END
 END vss.gds1619
 PIN vss.gds1620
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.242 15.695 71.282 15.895 ;
 END
 END vss.gds1620
 PIN vss.gds1621
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.57 15.695 70.61 15.895 ;
 END
 END vss.gds1621
 PIN vss.gds1622
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 18.1735 71.43 18.3735 ;
 END
 END vss.gds1622
 PIN vss.gds1623
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 18.1735 72.102 18.3735 ;
 END
 END vss.gds1623
 PIN vss.gds1624
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 18.1735 72.774 18.3735 ;
 END
 END vss.gds1624
 PIN vss.gds1625
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 18.1735 70.758 18.3735 ;
 END
 END vss.gds1625
 PIN vss.gds1626
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 18.1735 74.118 18.3735 ;
 END
 END vss.gds1626
 PIN vss.gds1627
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 18.1735 74.79 18.3735 ;
 END
 END vss.gds1627
 PIN vss.gds1628
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 18.1735 73.446 18.3735 ;
 END
 END vss.gds1628
 PIN vss.gds1629
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 74.564 18.493 74.62 18.693 ;
 RECT 74.06 18.483 74.116 18.683 ;
 RECT 73.892 18.493 73.948 18.693 ;
 RECT 73.388 18.483 73.444 18.683 ;
 RECT 73.22 18.493 73.276 18.693 ;
 RECT 72.716 18.483 72.772 18.683 ;
 RECT 72.548 18.493 72.604 18.693 ;
 RECT 72.044 18.483 72.1 18.683 ;
 RECT 71.876 18.493 71.932 18.693 ;
 RECT 71.372 18.483 71.428 18.683 ;
 RECT 71.204 18.493 71.26 18.693 ;
 RECT 70.7 18.483 70.756 18.683 ;
 RECT 70.532 18.493 70.588 18.693 ;
 RECT 74.396 15.721 74.452 15.921 ;
 RECT 74.228 15.721 74.284 15.921 ;
 RECT 74.564 15.736 74.62 15.936 ;
 RECT 73.724 15.721 73.78 15.921 ;
 RECT 73.556 15.721 73.612 15.921 ;
 RECT 73.892 15.736 73.948 15.936 ;
 RECT 74.06 15.736 74.116 15.936 ;
 RECT 73.052 15.721 73.108 15.921 ;
 RECT 72.884 15.721 72.94 15.921 ;
 RECT 73.22 15.736 73.276 15.936 ;
 RECT 73.388 15.736 73.444 15.936 ;
 RECT 72.38 15.721 72.436 15.921 ;
 RECT 72.212 15.721 72.268 15.921 ;
 RECT 72.548 15.736 72.604 15.936 ;
 RECT 72.716 15.736 72.772 15.936 ;
 RECT 71.708 15.721 71.764 15.921 ;
 RECT 71.54 15.721 71.596 15.921 ;
 RECT 71.876 15.736 71.932 15.936 ;
 RECT 72.044 15.736 72.1 15.936 ;
 RECT 71.036 15.721 71.092 15.921 ;
 RECT 70.868 15.721 70.924 15.921 ;
 RECT 71.204 15.736 71.26 15.936 ;
 RECT 71.372 15.736 71.428 15.936 ;
 RECT 70.364 15.721 70.42 15.921 ;
 RECT 70.532 15.736 70.588 15.936 ;
 RECT 70.7 15.736 70.756 15.936 ;
 RECT 74.396 16.795 74.452 16.995 ;
 RECT 74.228 16.795 74.284 16.995 ;
 RECT 74.732 15.736 74.788 15.936 ;
 RECT 74.732 18.483 74.788 18.683 ;
 RECT 74.732 16.795 74.788 16.995 ;
 RECT 74.564 16.795 74.62 16.995 ;
 RECT 73.724 16.795 73.78 16.995 ;
 RECT 73.556 16.795 73.612 16.995 ;
 RECT 74.06 16.795 74.116 16.995 ;
 RECT 73.892 16.795 73.948 16.995 ;
 RECT 73.052 16.795 73.108 16.995 ;
 RECT 72.884 16.795 72.94 16.995 ;
 RECT 73.388 16.795 73.444 16.995 ;
 RECT 73.22 16.795 73.276 16.995 ;
 RECT 72.38 16.795 72.436 16.995 ;
 RECT 72.212 16.795 72.268 16.995 ;
 RECT 72.716 16.795 72.772 16.995 ;
 RECT 72.548 16.795 72.604 16.995 ;
 RECT 71.708 16.795 71.764 16.995 ;
 RECT 71.54 16.795 71.596 16.995 ;
 RECT 72.044 16.795 72.1 16.995 ;
 RECT 71.876 16.795 71.932 16.995 ;
 RECT 71.036 16.795 71.092 16.995 ;
 RECT 70.868 16.795 70.924 16.995 ;
 RECT 71.372 16.795 71.428 16.995 ;
 RECT 71.204 16.795 71.26 16.995 ;
 RECT 70.364 16.795 70.42 16.995 ;
 RECT 70.7 16.795 70.756 16.995 ;
 RECT 70.532 16.795 70.588 16.995 ;
 END
 END vss.gds1629
 PIN vss.gds1630
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 23.469 0.29 23.669 ;
 END
 END vss.gds1630
 PIN vss.gds1631
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 25.357 2.962 25.557 ;
 END
 END vss.gds1631
 PIN vss.gds1632
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 21.577 2.962 21.777 ;
 END
 END vss.gds1632
 PIN vss.gds1633
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 24.097 2.962 24.297 ;
 END
 END vss.gds1633
 PIN vss.gds1634
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 23.696 3.142 23.896 ;
 END
 END vss.gds1634
 PIN vss.gds1635
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 22.436 3.142 22.636 ;
 END
 END vss.gds1635
 PIN vss.gds1636
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 24.956 3.142 25.156 ;
 END
 END vss.gds1636
 PIN vss.gds1637
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 22.837 2.962 23.037 ;
 END
 END vss.gds1637
 PIN vss.gds1638
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.286 20.947 3.326 21.147 ;
 END
 END vss.gds1638
 PIN vss.gds1639
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 21.176 3.142 21.376 ;
 END
 END vss.gds1639
 PIN vss.gds1640
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.442 20.541 4.482 20.741 ;
 END
 END vss.gds1640
 PIN vss.gds1641
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.414 21.223 3.454 21.423 ;
 END
 END vss.gds1641
 PIN vss.gds1642
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 23.262 0.602 23.462 ;
 END
 END vss.gds1642
 PIN vss.gds1643
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 23.061 0.942 23.261 ;
 END
 END vss.gds1643
 PIN vss.gds1644
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 23.605 1.282 23.805 ;
 END
 END vss.gds1644
 PIN vss.gds1645
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 23.4905 2.122 23.6905 ;
 END
 END vss.gds1645
 PIN vss.gds1646
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.754 23.467 3.794 23.667 ;
 END
 END vss.gds1646
 PIN vss.gds1647
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 23.467 5.074 23.667 ;
 END
 END vss.gds1647
 PIN vss.gds1648
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 23.467 4.194 23.667 ;
 END
 END vss.gds1648
 PIN vss.gds1649
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.57 20.744 4.61 20.944 ;
 END
 END vss.gds1649
 PIN vss.gds1650
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 23.3635 4.002 23.5635 ;
 END
 END vss.gds1650
 PIN vss.gds1651
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 23.3635 5.282 23.5635 ;
 END
 END vss.gds1651
 PIN vss.gds1652
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.562 20.6445 3.602 20.8445 ;
 END
 END vss.gds1652
 PIN vss.gds1653
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 22.772 2.302 22.972 ;
 END
 END vss.gds1653
 PIN vss.gds1654
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 23.5245 1.462 23.7245 ;
 END
 END vss.gds1654
 PIN vss.gds1655
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 23.1615 0.718 23.3615 ;
 END
 END vss.gds1655
 PIN vss.gds1656
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 2.576 21.5775 2.632 21.7775 ;
 RECT 2.408 21.5775 2.464 21.7775 ;
 RECT 2.996 21.5775 3.052 21.7775 ;
 RECT 3.332 21.669 3.388 21.869 ;
 RECT 3.5 21.6255 3.556 21.8255 ;
 RECT 0.98 21.4925 1.036 21.6925 ;
 RECT 2.072 21.493 2.128 21.693 ;
 RECT 2.576 22.8375 2.632 23.0375 ;
 RECT 2.408 22.8375 2.464 23.0375 ;
 RECT 2.996 22.8375 3.052 23.0375 ;
 RECT 3.332 22.929 3.388 23.129 ;
 RECT 3.5 22.8855 3.556 23.0855 ;
 RECT 0.98 22.7525 1.036 22.9525 ;
 RECT 2.072 22.753 2.128 22.953 ;
 RECT 2.576 24.0975 2.632 24.2975 ;
 RECT 2.408 24.0975 2.464 24.2975 ;
 RECT 2.996 24.0975 3.052 24.2975 ;
 RECT 3.332 24.189 3.388 24.389 ;
 RECT 3.5 24.1455 3.556 24.3455 ;
 RECT 0.98 24.0125 1.036 24.2125 ;
 RECT 2.072 24.013 2.128 24.213 ;
 RECT 2.576 25.3575 2.632 25.5575 ;
 RECT 2.408 25.3575 2.464 25.5575 ;
 RECT 2.996 25.3575 3.052 25.5575 ;
 RECT 3.5 25.4055 3.556 25.6055 ;
 RECT 0.98 25.2725 1.036 25.4725 ;
 RECT 2.072 25.273 2.128 25.473 ;
 RECT 0.392 25.363 0.448 25.563 ;
 RECT 0.644 25.363 0.7 25.563 ;
 RECT 1.232 25.363 1.288 25.563 ;
 RECT 1.4 25.363 1.456 25.563 ;
 RECT 1.568 25.363 1.624 25.563 ;
 RECT 1.82 25.363 1.876 25.563 ;
 RECT 2.24 25.363 2.296 25.563 ;
 RECT 2.744 25.273 2.8 25.473 ;
 RECT 3.164 25.363 3.22 25.563 ;
 RECT 3.92 25.363 3.976 25.563 ;
 RECT 0.392 24.103 0.448 24.303 ;
 RECT 0.812 24.189 0.868 24.389 ;
 RECT 0.644 24.103 0.7 24.303 ;
 RECT 1.232 24.103 1.288 24.303 ;
 RECT 1.4 24.103 1.456 24.303 ;
 RECT 1.568 24.103 1.624 24.303 ;
 RECT 1.82 24.103 1.876 24.303 ;
 RECT 2.24 24.103 2.296 24.303 ;
 RECT 2.744 24.013 2.8 24.213 ;
 RECT 3.164 24.103 3.22 24.303 ;
 RECT 3.92 24.103 3.976 24.303 ;
 RECT 3.752 24.373 3.808 24.573 ;
 RECT 4.508 24.3025 4.564 24.5025 ;
 RECT 0.392 22.843 0.448 23.043 ;
 RECT 0.812 22.929 0.868 23.129 ;
 RECT 0.644 22.843 0.7 23.043 ;
 RECT 1.232 22.843 1.288 23.043 ;
 RECT 1.4 22.843 1.456 23.043 ;
 RECT 1.568 22.843 1.624 23.043 ;
 RECT 1.82 22.843 1.876 23.043 ;
 RECT 2.24 22.843 2.296 23.043 ;
 RECT 2.744 22.753 2.8 22.953 ;
 RECT 3.164 22.843 3.22 23.043 ;
 RECT 3.92 22.843 3.976 23.043 ;
 RECT 3.752 23.113 3.808 23.313 ;
 RECT 4.508 23.0425 4.564 23.2425 ;
 RECT 0.392 21.583 0.448 21.783 ;
 RECT 0.812 21.669 0.868 21.869 ;
 RECT 0.644 21.583 0.7 21.783 ;
 RECT 1.232 21.583 1.288 21.783 ;
 RECT 1.4 21.583 1.456 21.783 ;
 RECT 1.568 21.583 1.624 21.783 ;
 RECT 1.82 21.583 1.876 21.783 ;
 RECT 2.24 21.583 2.296 21.783 ;
 RECT 2.744 21.493 2.8 21.693 ;
 RECT 3.164 21.583 3.22 21.783 ;
 RECT 3.92 21.583 3.976 21.783 ;
 RECT 3.752 21.853 3.808 22.053 ;
 RECT 4.508 21.7825 4.564 21.9825 ;
 RECT 3.752 20.593 3.808 20.793 ;
 RECT 4.508 20.5225 4.564 20.7225 ;
 END
 END vss.gds1656
 PIN vss.gds1657
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.134 21.1635 10.194 21.3635 ;
 END
 END vss.gds1657
 PIN vss.gds1658
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.966 21.1635 10.026 21.3635 ;
 END
 END vss.gds1658
 PIN vss.gds1659
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.798 21.1635 9.858 21.3635 ;
 END
 END vss.gds1659
 PIN vss.gds1660
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.462 21.1635 9.522 21.3635 ;
 END
 END vss.gds1660
 PIN vss.gds1661
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.294 21.1635 9.354 21.3635 ;
 END
 END vss.gds1661
 PIN vss.gds1662
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.79 21.1635 8.85 21.3635 ;
 END
 END vss.gds1662
 PIN vss.gds1663
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.622 21.1635 8.682 21.3635 ;
 END
 END vss.gds1663
 PIN vss.gds1664
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.454 21.1635 8.514 21.3635 ;
 END
 END vss.gds1664
 PIN vss.gds1665
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.118 21.1635 8.178 21.3635 ;
 END
 END vss.gds1665
 PIN vss.gds1666
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.95 21.1635 8.01 21.3635 ;
 END
 END vss.gds1666
 PIN vss.gds1667
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.782 21.1635 7.842 21.3635 ;
 END
 END vss.gds1667
 PIN vss.gds1668
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.126 21.1635 9.186 21.3635 ;
 END
 END vss.gds1668
 PIN vss.gds1669
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.446 21.1635 7.506 21.3635 ;
 END
 END vss.gds1669
 PIN vss.gds1670
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.278 21.1635 7.338 21.3635 ;
 END
 END vss.gds1670
 PIN vss.gds1671
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 22.9275 9.69 23.1275 ;
 END
 END vss.gds1671
 PIN vss.gds1672
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 22.9275 8.346 23.1275 ;
 END
 END vss.gds1672
 PIN vss.gds1673
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 22.9275 9.018 23.1275 ;
 END
 END vss.gds1673
 PIN vss.gds1674
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 22.9275 7.674 23.1275 ;
 END
 END vss.gds1674
 PIN vss.gds1675
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.11 21.1635 7.17 21.3635 ;
 END
 END vss.gds1675
 PIN vss.gds1676
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 23.467 5.474 23.667 ;
 END
 END vss.gds1676
 PIN vss.gds1677
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 23.467 5.986 23.667 ;
 END
 END vss.gds1677
 PIN vss.gds1678
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 23.264 6.178 23.464 ;
 END
 END vss.gds1678
 PIN vss.gds1679
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 23.467 5.73 23.667 ;
 END
 END vss.gds1679
 PIN vss.gds1680
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 23.263 6.434 23.463 ;
 END
 END vss.gds1680
 PIN vss.gds1681
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 6.524 25.325 6.58 25.525 ;
 RECT 6.524 24.065 6.58 24.265 ;
 RECT 6.524 22.805 6.58 23.005 ;
 RECT 6.524 21.545 6.58 21.745 ;
 RECT 6.692 20.608 6.748 20.808 ;
 RECT 6.692 21.868 6.748 22.068 ;
 RECT 6.692 23.128 6.748 23.328 ;
 RECT 6.692 24.388 6.748 24.588 ;
 RECT 6.608 24.373 6.664 24.573 ;
 RECT 6.608 23.113 6.664 23.313 ;
 RECT 6.608 21.853 6.664 22.053 ;
 RECT 6.608 20.593 6.664 20.793 ;
 END
 END vss.gds1681
 PIN vss.gds1682
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 22.082 13.898 22.282 ;
 END
 END vss.gds1682
 PIN vss.gds1683
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 22.122 14.87 22.322 ;
 END
 END vss.gds1683
 PIN vss.gds1684
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 20.822 13.898 21.022 ;
 END
 END vss.gds1684
 PIN vss.gds1685
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 20.862 14.87 21.062 ;
 END
 END vss.gds1685
 PIN vss.gds1686
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 24.602 13.898 24.802 ;
 END
 END vss.gds1686
 PIN vss.gds1687
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 24.642 14.87 24.842 ;
 END
 END vss.gds1687
 PIN vss.gds1688
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 23.342 13.898 23.542 ;
 END
 END vss.gds1688
 PIN vss.gds1689
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 23.382 14.87 23.582 ;
 END
 END vss.gds1689
 PIN vss.gds1690
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.15 21.1635 12.21 21.3635 ;
 END
 END vss.gds1690
 PIN vss.gds1691
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.982 21.1635 12.042 21.3635 ;
 END
 END vss.gds1691
 PIN vss.gds1692
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.814 21.1635 11.874 21.3635 ;
 END
 END vss.gds1692
 PIN vss.gds1693
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.478 21.1635 11.538 21.3635 ;
 END
 END vss.gds1693
 PIN vss.gds1694
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.31 21.1635 11.37 21.3635 ;
 END
 END vss.gds1694
 PIN vss.gds1695
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.142 21.1635 11.202 21.3635 ;
 END
 END vss.gds1695
 PIN vss.gds1696
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.806 21.1635 10.866 21.3635 ;
 END
 END vss.gds1696
 PIN vss.gds1697
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.638 21.1635 10.698 21.3635 ;
 END
 END vss.gds1697
 PIN vss.gds1698
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.47 21.1635 10.53 21.3635 ;
 END
 END vss.gds1698
 PIN vss.gds1699
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 22.9275 13.658 23.1275 ;
 END
 END vss.gds1699
 PIN vss.gds1700
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 21.8495 13.058 22.0495 ;
 END
 END vss.gds1700
 PIN vss.gds1701
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.262 24.156 13.318 24.356 ;
 END
 END vss.gds1701
 PIN vss.gds1702
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 22.9275 11.706 23.1275 ;
 END
 END vss.gds1702
 PIN vss.gds1703
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 22.9275 11.034 23.1275 ;
 END
 END vss.gds1703
 PIN vss.gds1704
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 23.22 15.162 23.42 ;
 END
 END vss.gds1704
 PIN vss.gds1705
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 22.9275 10.362 23.1275 ;
 END
 END vss.gds1705
 PIN vss.gds1706
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 23.22 14.498 23.42 ;
 END
 END vss.gds1706
 PIN vss.gds1707
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 23.0835 12.818 23.2835 ;
 END
 END vss.gds1707
 PIN vss.gds1708
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 22.765 12.378 22.965 ;
 END
 END vss.gds1708
 PIN vss.gds1709
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 23.467 12.59 23.667 ;
 END
 END vss.gds1709
 PIN vss.gds1710
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 14 22.26 14.056 22.433 ;
 RECT 14.168 22.233 14.224 22.433 ;
 RECT 14 23.52 14.056 23.693 ;
 RECT 14.168 23.493 14.224 23.693 ;
 RECT 14 24.78 14.056 24.953 ;
 RECT 14.168 24.753 14.224 24.953 ;
 RECT 14.336 21.593 14.392 21.793 ;
 RECT 14.168 21.593 14.224 21.793 ;
 RECT 14.336 25.373 14.392 25.573 ;
 RECT 14.168 25.373 14.224 25.573 ;
 RECT 14.336 24.113 14.392 24.313 ;
 RECT 14.168 24.113 14.224 24.313 ;
 RECT 14.336 22.853 14.392 23.053 ;
 RECT 14.168 22.853 14.224 23.053 ;
 RECT 15.008 24.323 15.064 24.523 ;
 RECT 14.84 24.797 14.896 24.962 ;
 RECT 14.672 24.797 14.728 24.962 ;
 RECT 13.664 24.247 13.72 24.447 ;
 RECT 13.664 22.987 13.72 23.187 ;
 RECT 15.008 23.063 15.064 23.263 ;
 RECT 14.84 23.537 14.896 23.702 ;
 RECT 14.672 23.537 14.728 23.702 ;
 RECT 14 21 14.056 21.173 ;
 RECT 14.168 20.973 14.224 21.173 ;
 RECT 14.84 21.017 14.896 21.182 ;
 RECT 14.672 21.017 14.728 21.182 ;
 RECT 15.008 20.543 15.064 20.743 ;
 RECT 13.664 20.467 13.72 20.667 ;
 RECT 15.008 21.803 15.064 22.003 ;
 RECT 14.84 22.277 14.896 22.442 ;
 RECT 14.672 22.277 14.728 22.442 ;
 RECT 13.664 21.727 13.72 21.927 ;
 RECT 15.176 21.2435 15.232 21.4435 ;
 RECT 12.824 21.028 12.88 21.228 ;
 RECT 13.496 21.039 13.552 21.239 ;
 RECT 13.328 20.977 13.384 21.177 ;
 RECT 13.16 21.028 13.216 21.228 ;
 RECT 12.488 21.058 12.544 21.258 ;
 RECT 12.992 21.028 13.048 21.228 ;
 RECT 12.656 21.058 12.712 21.258 ;
 END
 END vss.gds1710
 PIN vss.gds1711
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.986 20.947 18.026 21.147 ;
 END
 END vss.gds1711
 PIN vss.gds1712
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 22.837 16.146 23.037 ;
 END
 END vss.gds1712
 PIN vss.gds1713
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 24.84 15.418 25.04 ;
 END
 END vss.gds1713
 PIN vss.gds1714
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 24.097 16.146 24.297 ;
 END
 END vss.gds1714
 PIN vss.gds1715
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.438 23.7395 17.494 23.9395 ;
 END
 END vss.gds1715
 PIN vss.gds1716
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.038 21.1635 19.098 21.3635 ;
 END
 END vss.gds1716
 PIN vss.gds1717
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.206 21.1635 19.266 21.3635 ;
 END
 END vss.gds1717
 PIN vss.gds1718
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.374 21.1635 19.434 21.3635 ;
 END
 END vss.gds1718
 PIN vss.gds1719
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 22.9275 20.274 23.1275 ;
 END
 END vss.gds1719
 PIN vss.gds1720
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 25.357 16.146 25.557 ;
 END
 END vss.gds1720
 PIN vss.gds1721
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.702 21.1635 18.762 21.3635 ;
 END
 END vss.gds1721
 PIN vss.gds1722
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.71 21.1635 19.77 21.3635 ;
 END
 END vss.gds1722
 PIN vss.gds1723
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.878 21.1635 19.938 21.3635 ;
 END
 END vss.gds1723
 PIN vss.gds1724
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.534 21.1635 18.594 21.3635 ;
 END
 END vss.gds1724
 PIN vss.gds1725
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 21.636 16.814 21.836 ;
 END
 END vss.gds1725
 PIN vss.gds1726
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 24.8475 17.314 25.0475 ;
 END
 END vss.gds1726
 PIN vss.gds1727
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.366 21.1635 18.426 21.3635 ;
 END
 END vss.gds1727
 PIN vss.gds1728
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.046 21.1635 20.106 21.3635 ;
 END
 END vss.gds1728
 PIN vss.gds1729
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 21.577 16.146 21.777 ;
 END
 END vss.gds1729
 PIN vss.gds1730
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 22.9275 19.602 23.1275 ;
 END
 END vss.gds1730
 PIN vss.gds1731
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 22.9275 18.93 23.1275 ;
 END
 END vss.gds1731
 PIN vss.gds1732
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 22.8865 16.994 23.0865 ;
 END
 END vss.gds1732
 PIN vss.gds1733
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 23.22 15.842 23.42 ;
 END
 END vss.gds1733
 PIN vss.gds1734
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 23.0835 17.834 23.2835 ;
 END
 END vss.gds1734
 PIN vss.gds1735
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 23.4905 16.49 23.6905 ;
 END
 END vss.gds1735
 PIN vss.gds1736
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 22.765 18.258 22.965 ;
 END
 END vss.gds1736
 PIN vss.gds1737
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 15.596 25.024 15.652 25.224 ;
 RECT 15.848 25.027 15.904 25.227 ;
 RECT 15.596 21.244 15.652 21.444 ;
 RECT 15.848 21.247 15.904 21.447 ;
 RECT 16.52 22.28 16.576 22.433 ;
 RECT 15.764 22.277 15.82 22.442 ;
 RECT 15.596 22.277 15.652 22.442 ;
 RECT 15.596 22.504 15.652 22.704 ;
 RECT 15.848 22.507 15.904 22.707 ;
 RECT 16.52 23.54 16.576 23.693 ;
 RECT 15.764 23.537 15.82 23.702 ;
 RECT 15.596 23.537 15.652 23.702 ;
 RECT 15.596 23.764 15.652 23.964 ;
 RECT 15.848 23.767 15.904 23.967 ;
 RECT 16.52 24.8 16.576 24.953 ;
 RECT 15.764 24.797 15.82 24.962 ;
 RECT 15.596 24.797 15.652 24.962 ;
 RECT 16.352 23.1635 16.408 23.3635 ;
 RECT 16.856 22.9115 16.912 23.1115 ;
 RECT 15.428 24.323 15.484 24.523 ;
 RECT 16.352 24.4235 16.408 24.6235 ;
 RECT 16.856 24.1715 16.912 24.3715 ;
 RECT 15.428 23.063 15.484 23.263 ;
 RECT 16.52 21.02 16.576 21.173 ;
 RECT 15.764 21.017 15.82 21.182 ;
 RECT 15.596 21.017 15.652 21.182 ;
 RECT 15.428 20.543 15.484 20.743 ;
 RECT 16.352 20.6435 16.408 20.8435 ;
 RECT 15.428 21.803 15.484 22.003 ;
 RECT 16.352 21.9035 16.408 22.1035 ;
 RECT 16.856 21.6515 16.912 21.8515 ;
 RECT 16.856 25.4315 16.912 25.6315 ;
 RECT 17.864 21.058 17.92 21.258 ;
 RECT 17.696 21.0655 17.752 21.2655 ;
 RECT 17.528 21.058 17.584 21.258 ;
 RECT 17.36 21.058 17.416 21.258 ;
 RECT 17.192 21.058 17.248 21.258 ;
 RECT 18.032 21.058 18.088 21.258 ;
 RECT 17.024 21.173 17.08 21.373 ;
 END
 END vss.gds1737
 PIN vss.gds1738
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.17 21.1635 25.23 21.3635 ;
 END
 END vss.gds1738
 PIN vss.gds1739
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.002 21.1635 25.062 21.3635 ;
 END
 END vss.gds1739
 PIN vss.gds1740
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.834 21.1635 24.894 21.3635 ;
 END
 END vss.gds1740
 PIN vss.gds1741
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.498 21.1635 24.558 21.3635 ;
 END
 END vss.gds1741
 PIN vss.gds1742
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.33 21.1635 24.39 21.3635 ;
 END
 END vss.gds1742
 PIN vss.gds1743
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.162 21.1635 24.222 21.3635 ;
 END
 END vss.gds1743
 PIN vss.gds1744
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.382 21.1635 20.442 21.3635 ;
 END
 END vss.gds1744
 PIN vss.gds1745
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.55 21.1635 20.61 21.3635 ;
 END
 END vss.gds1745
 PIN vss.gds1746
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.718 21.1635 20.778 21.3635 ;
 END
 END vss.gds1746
 PIN vss.gds1747
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.054 21.1635 21.114 21.3635 ;
 END
 END vss.gds1747
 PIN vss.gds1748
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.222 21.1635 21.282 21.3635 ;
 END
 END vss.gds1748
 PIN vss.gds1749
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.39 21.1635 21.45 21.3635 ;
 END
 END vss.gds1749
 PIN vss.gds1750
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.726 21.1635 21.786 21.3635 ;
 END
 END vss.gds1750
 PIN vss.gds1751
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.894 21.1635 21.954 21.3635 ;
 END
 END vss.gds1751
 PIN vss.gds1752
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.062 21.1635 22.122 21.3635 ;
 END
 END vss.gds1752
 PIN vss.gds1753
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.398 21.1635 22.458 21.3635 ;
 END
 END vss.gds1753
 PIN vss.gds1754
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.566 21.1635 22.626 21.3635 ;
 END
 END vss.gds1754
 PIN vss.gds1755
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.734 21.1635 22.794 21.3635 ;
 END
 END vss.gds1755
 PIN vss.gds1756
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.07 21.1635 23.13 21.3635 ;
 END
 END vss.gds1756
 PIN vss.gds1757
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.238 21.1635 23.298 21.3635 ;
 END
 END vss.gds1757
 PIN vss.gds1758
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.406 21.1635 23.466 21.3635 ;
 END
 END vss.gds1758
 PIN vss.gds1759
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 22.9275 24.726 23.1275 ;
 END
 END vss.gds1759
 PIN vss.gds1760
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 22.9275 22.962 23.1275 ;
 END
 END vss.gds1760
 PIN vss.gds1761
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 22.9275 22.29 23.1275 ;
 END
 END vss.gds1761
 PIN vss.gds1762
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 22.9275 21.618 23.1275 ;
 END
 END vss.gds1762
 PIN vss.gds1763
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 22.9275 20.946 23.1275 ;
 END
 END vss.gds1763
 PIN vss.gds1764
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 22.9275 23.634 23.1275 ;
 END
 END vss.gds1764
 PIN vss.gds1765
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 23.912 23 23.968 23.2 ;
 RECT 23.912 24.26 23.968 24.46 ;
 RECT 23.912 20.48 23.968 20.68 ;
 RECT 23.912 21.74 23.968 21.94 ;
 RECT 23.744 23.07 23.8 23.27 ;
 END
 END vss.gds1765
 PIN vss.gds1766
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.202 21.1635 29.262 21.3635 ;
 END
 END vss.gds1766
 PIN vss.gds1767
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.034 21.1635 29.094 21.3635 ;
 END
 END vss.gds1767
 PIN vss.gds1768
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.866 21.1635 28.926 21.3635 ;
 END
 END vss.gds1768
 PIN vss.gds1769
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.53 21.1635 28.59 21.3635 ;
 END
 END vss.gds1769
 PIN vss.gds1770
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.362 21.1635 28.422 21.3635 ;
 END
 END vss.gds1770
 PIN vss.gds1771
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.194 21.1635 28.254 21.3635 ;
 END
 END vss.gds1771
 PIN vss.gds1772
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.858 21.1635 27.918 21.3635 ;
 END
 END vss.gds1772
 PIN vss.gds1773
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.69 21.1635 27.75 21.3635 ;
 END
 END vss.gds1773
 PIN vss.gds1774
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.522 21.1635 27.582 21.3635 ;
 END
 END vss.gds1774
 PIN vss.gds1775
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.186 21.1635 27.246 21.3635 ;
 END
 END vss.gds1775
 PIN vss.gds1776
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.018 21.1635 27.078 21.3635 ;
 END
 END vss.gds1776
 PIN vss.gds1777
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.85 21.1635 26.91 21.3635 ;
 END
 END vss.gds1777
 PIN vss.gds1778
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.514 21.1635 26.574 21.3635 ;
 END
 END vss.gds1778
 PIN vss.gds1779
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.346 21.1635 26.406 21.3635 ;
 END
 END vss.gds1779
 PIN vss.gds1780
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.178 21.1635 26.238 21.3635 ;
 END
 END vss.gds1780
 PIN vss.gds1781
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.842 21.1635 25.902 21.3635 ;
 END
 END vss.gds1781
 PIN vss.gds1782
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.674 21.1635 25.734 21.3635 ;
 END
 END vss.gds1782
 PIN vss.gds1783
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.506 21.1635 25.566 21.3635 ;
 END
 END vss.gds1783
 PIN vss.gds1784
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 22.765 29.43 22.965 ;
 END
 END vss.gds1784
 PIN vss.gds1785
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 22.9275 28.758 23.1275 ;
 END
 END vss.gds1785
 PIN vss.gds1786
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 22.9275 28.086 23.1275 ;
 END
 END vss.gds1786
 PIN vss.gds1787
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 22.9275 27.414 23.1275 ;
 END
 END vss.gds1787
 PIN vss.gds1788
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 22.9275 26.742 23.1275 ;
 END
 END vss.gds1788
 PIN vss.gds1789
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 22.9275 26.07 23.1275 ;
 END
 END vss.gds1789
 PIN vss.gds1790
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 22.9275 25.398 23.1275 ;
 END
 END vss.gds1790
 PIN vss.gds1791
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 21.8495 30.11 22.0495 ;
 END
 END vss.gds1791
 PIN vss.gds1792
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 23.0835 29.87 23.2835 ;
 END
 END vss.gds1792
 PIN vss.gds1793
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 23.467 29.642 23.667 ;
 END
 END vss.gds1793
 PIN vss.gds1794
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.876 21.028 29.932 21.228 ;
 RECT 30.212 21.028 30.268 21.228 ;
 RECT 29.54 21.058 29.596 21.258 ;
 RECT 29.708 21.058 29.764 21.258 ;
 RECT 30.044 21.028 30.1 21.228 ;
 END
 END vss.gds1794
 PIN vss.gds1795
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 22.122 31.922 22.322 ;
 END
 END vss.gds1795
 PIN vss.gds1796
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 20.822 30.95 21.022 ;
 END
 END vss.gds1796
 PIN vss.gds1797
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 20.862 31.922 21.062 ;
 END
 END vss.gds1797
 PIN vss.gds1798
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 24.642 31.922 24.842 ;
 END
 END vss.gds1798
 PIN vss.gds1799
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 23.342 30.95 23.542 ;
 END
 END vss.gds1799
 PIN vss.gds1800
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 23.382 31.922 23.582 ;
 END
 END vss.gds1800
 PIN vss.gds1801
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 24.84 32.47 25.04 ;
 END
 END vss.gds1801
 PIN vss.gds1802
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 24.602 30.95 24.802 ;
 END
 END vss.gds1802
 PIN vss.gds1803
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 24.097 33.198 24.297 ;
 END
 END vss.gds1803
 PIN vss.gds1804
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 22.837 33.198 23.037 ;
 END
 END vss.gds1804
 PIN vss.gds1805
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.038 20.947 35.078 21.147 ;
 END
 END vss.gds1805
 PIN vss.gds1806
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.314 24.156 30.37 24.356 ;
 END
 END vss.gds1806
 PIN vss.gds1807
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 23.22 32.894 23.42 ;
 END
 END vss.gds1807
 PIN vss.gds1808
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 23.22 32.214 23.42 ;
 END
 END vss.gds1808
 PIN vss.gds1809
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.49 23.7395 34.546 23.9395 ;
 END
 END vss.gds1809
 PIN vss.gds1810
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 22.9275 30.71 23.1275 ;
 END
 END vss.gds1810
 PIN vss.gds1811
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 21.636 33.866 21.836 ;
 END
 END vss.gds1811
 PIN vss.gds1812
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 21.577 33.198 21.777 ;
 END
 END vss.gds1812
 PIN vss.gds1813
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 25.357 33.198 25.557 ;
 END
 END vss.gds1813
 PIN vss.gds1814
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 23.4905 33.542 23.6905 ;
 END
 END vss.gds1814
 PIN vss.gds1815
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 24.8475 34.366 25.0475 ;
 END
 END vss.gds1815
 PIN vss.gds1816
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 22.082 30.95 22.282 ;
 END
 END vss.gds1816
 PIN vss.gds1817
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 23.22 31.55 23.42 ;
 END
 END vss.gds1817
 PIN vss.gds1818
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 23.0835 34.886 23.2835 ;
 END
 END vss.gds1818
 PIN vss.gds1819
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 22.8865 34.046 23.0865 ;
 END
 END vss.gds1819
 PIN vss.gds1820
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 32.648 25.024 32.704 25.224 ;
 RECT 32.9 25.027 32.956 25.227 ;
 RECT 32.648 21.244 32.704 21.444 ;
 RECT 32.9 21.247 32.956 21.447 ;
 RECT 33.572 22.28 33.628 22.433 ;
 RECT 31.052 22.26 31.108 22.433 ;
 RECT 31.22 22.233 31.276 22.433 ;
 RECT 32.816 22.277 32.872 22.442 ;
 RECT 32.648 22.277 32.704 22.442 ;
 RECT 31.892 22.277 31.948 22.442 ;
 RECT 31.724 22.277 31.78 22.442 ;
 RECT 33.572 21.02 33.628 21.173 ;
 RECT 31.052 21 31.108 21.173 ;
 RECT 31.22 20.973 31.276 21.173 ;
 RECT 32.816 21.017 32.872 21.182 ;
 RECT 32.648 21.017 32.704 21.182 ;
 RECT 31.892 21.017 31.948 21.182 ;
 RECT 31.724 21.017 31.78 21.182 ;
 RECT 33.572 23.54 33.628 23.693 ;
 RECT 31.052 23.52 31.108 23.693 ;
 RECT 31.22 23.493 31.276 23.693 ;
 RECT 32.816 23.537 32.872 23.702 ;
 RECT 32.648 23.537 32.704 23.702 ;
 RECT 31.892 23.537 31.948 23.702 ;
 RECT 31.724 23.537 31.78 23.702 ;
 RECT 32.648 23.764 32.704 23.964 ;
 RECT 32.9 23.767 32.956 23.967 ;
 RECT 33.572 24.8 33.628 24.953 ;
 RECT 31.052 24.78 31.108 24.953 ;
 RECT 31.22 24.753 31.276 24.953 ;
 RECT 32.816 24.797 32.872 24.962 ;
 RECT 32.648 24.797 32.704 24.962 ;
 RECT 31.892 24.797 31.948 24.962 ;
 RECT 31.724 24.797 31.78 24.962 ;
 RECT 32.648 22.504 32.704 22.704 ;
 RECT 32.9 22.507 32.956 22.707 ;
 RECT 32.06 24.323 32.116 24.523 ;
 RECT 31.388 24.113 31.444 24.313 ;
 RECT 31.22 24.113 31.276 24.313 ;
 RECT 32.48 24.323 32.536 24.523 ;
 RECT 33.404 23.1635 33.46 23.3635 ;
 RECT 33.908 22.9115 33.964 23.1115 ;
 RECT 31.388 22.853 31.444 23.053 ;
 RECT 31.22 22.853 31.276 23.053 ;
 RECT 31.388 21.593 31.444 21.793 ;
 RECT 31.22 21.593 31.276 21.793 ;
 RECT 32.06 21.803 32.116 22.003 ;
 RECT 32.48 21.803 32.536 22.003 ;
 RECT 33.908 25.4315 33.964 25.6315 ;
 RECT 31.388 25.373 31.444 25.573 ;
 RECT 31.22 25.373 31.276 25.573 ;
 RECT 30.716 22.987 30.772 23.187 ;
 RECT 32.06 23.063 32.116 23.263 ;
 RECT 32.48 23.063 32.536 23.263 ;
 RECT 32.06 20.543 32.116 20.743 ;
 RECT 32.48 20.543 32.536 20.743 ;
 RECT 30.716 20.467 30.772 20.667 ;
 RECT 30.716 24.247 30.772 24.447 ;
 RECT 33.404 24.4235 33.46 24.6235 ;
 RECT 33.908 24.1715 33.964 24.3715 ;
 RECT 30.716 21.727 30.772 21.927 ;
 RECT 33.404 21.9035 33.46 22.1035 ;
 RECT 33.908 21.6515 33.964 21.8515 ;
 RECT 30.548 21.039 30.604 21.239 ;
 RECT 33.404 20.6435 33.46 20.8435 ;
 RECT 32.228 21.2435 32.284 21.4435 ;
 RECT 30.38 20.977 30.436 21.177 ;
 RECT 34.916 21.058 34.972 21.258 ;
 RECT 34.748 21.0655 34.804 21.2655 ;
 RECT 34.58 21.058 34.636 21.258 ;
 RECT 34.412 21.058 34.468 21.258 ;
 RECT 34.244 21.058 34.3 21.258 ;
 RECT 35.084 21.058 35.14 21.258 ;
 RECT 34.076 21.173 34.132 21.373 ;
 END
 END vss.gds1820
 PIN vss.gds1821
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.122 21.1635 40.182 21.3635 ;
 END
 END vss.gds1821
 PIN vss.gds1822
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.754 21.1635 35.814 21.3635 ;
 END
 END vss.gds1822
 PIN vss.gds1823
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.09 21.1635 36.15 21.3635 ;
 END
 END vss.gds1823
 PIN vss.gds1824
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.258 21.1635 36.318 21.3635 ;
 END
 END vss.gds1824
 PIN vss.gds1825
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.426 21.1635 36.486 21.3635 ;
 END
 END vss.gds1825
 PIN vss.gds1826
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.762 21.1635 36.822 21.3635 ;
 END
 END vss.gds1826
 PIN vss.gds1827
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.93 21.1635 36.99 21.3635 ;
 END
 END vss.gds1827
 PIN vss.gds1828
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.098 21.1635 37.158 21.3635 ;
 END
 END vss.gds1828
 PIN vss.gds1829
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.434 21.1635 37.494 21.3635 ;
 END
 END vss.gds1829
 PIN vss.gds1830
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.602 21.1635 37.662 21.3635 ;
 END
 END vss.gds1830
 PIN vss.gds1831
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.77 21.1635 37.83 21.3635 ;
 END
 END vss.gds1831
 PIN vss.gds1832
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.106 21.1635 38.166 21.3635 ;
 END
 END vss.gds1832
 PIN vss.gds1833
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.274 21.1635 38.334 21.3635 ;
 END
 END vss.gds1833
 PIN vss.gds1834
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.442 21.1635 38.502 21.3635 ;
 END
 END vss.gds1834
 PIN vss.gds1835
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 22.9275 37.998 23.1275 ;
 END
 END vss.gds1835
 PIN vss.gds1836
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 22.9275 37.326 23.1275 ;
 END
 END vss.gds1836
 PIN vss.gds1837
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 22.9275 38.67 23.1275 ;
 END
 END vss.gds1837
 PIN vss.gds1838
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.778 21.1635 38.838 21.3635 ;
 END
 END vss.gds1838
 PIN vss.gds1839
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.946 21.1635 39.006 21.3635 ;
 END
 END vss.gds1839
 PIN vss.gds1840
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.114 21.1635 39.174 21.3635 ;
 END
 END vss.gds1840
 PIN vss.gds1841
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.45 21.1635 39.51 21.3635 ;
 END
 END vss.gds1841
 PIN vss.gds1842
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.618 21.1635 39.678 21.3635 ;
 END
 END vss.gds1842
 PIN vss.gds1843
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.786 21.1635 39.846 21.3635 ;
 END
 END vss.gds1843
 PIN vss.gds1844
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.586 21.1635 35.646 21.3635 ;
 END
 END vss.gds1844
 PIN vss.gds1845
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.418 21.1635 35.478 21.3635 ;
 END
 END vss.gds1845
 PIN vss.gds1846
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 22.9275 36.654 23.1275 ;
 END
 END vss.gds1846
 PIN vss.gds1847
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 22.9275 39.342 23.1275 ;
 END
 END vss.gds1847
 PIN vss.gds1848
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 22.9275 40.014 23.1275 ;
 END
 END vss.gds1848
 PIN vss.gds1849
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 22.765 35.31 22.965 ;
 END
 END vss.gds1849
 PIN vss.gds1850
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 22.9275 35.982 23.1275 ;
 END
 END vss.gds1850
 PIN vss.gds1851
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.91 21.1635 44.97 21.3635 ;
 END
 END vss.gds1851
 PIN vss.gds1852
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.742 21.1635 44.802 21.3635 ;
 END
 END vss.gds1852
 PIN vss.gds1853
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.574 21.1635 44.634 21.3635 ;
 END
 END vss.gds1853
 PIN vss.gds1854
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.238 21.1635 44.298 21.3635 ;
 END
 END vss.gds1854
 PIN vss.gds1855
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.07 21.1635 44.13 21.3635 ;
 END
 END vss.gds1855
 PIN vss.gds1856
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.902 21.1635 43.962 21.3635 ;
 END
 END vss.gds1856
 PIN vss.gds1857
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.566 21.1635 43.626 21.3635 ;
 END
 END vss.gds1857
 PIN vss.gds1858
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.398 21.1635 43.458 21.3635 ;
 END
 END vss.gds1858
 PIN vss.gds1859
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.23 21.1635 43.29 21.3635 ;
 END
 END vss.gds1859
 PIN vss.gds1860
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.894 21.1635 42.954 21.3635 ;
 END
 END vss.gds1860
 PIN vss.gds1861
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.726 21.1635 42.786 21.3635 ;
 END
 END vss.gds1861
 PIN vss.gds1862
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.558 21.1635 42.618 21.3635 ;
 END
 END vss.gds1862
 PIN vss.gds1863
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.222 21.1635 42.282 21.3635 ;
 END
 END vss.gds1863
 PIN vss.gds1864
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.054 21.1635 42.114 21.3635 ;
 END
 END vss.gds1864
 PIN vss.gds1865
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.886 21.1635 41.946 21.3635 ;
 END
 END vss.gds1865
 PIN vss.gds1866
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.55 21.1635 41.61 21.3635 ;
 END
 END vss.gds1866
 PIN vss.gds1867
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.382 21.1635 41.442 21.3635 ;
 END
 END vss.gds1867
 PIN vss.gds1868
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.214 21.1635 41.274 21.3635 ;
 END
 END vss.gds1868
 PIN vss.gds1869
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.29 21.1635 40.35 21.3635 ;
 END
 END vss.gds1869
 PIN vss.gds1870
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.458 21.1635 40.518 21.3635 ;
 END
 END vss.gds1870
 PIN vss.gds1871
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 22.9275 45.138 23.1275 ;
 END
 END vss.gds1871
 PIN vss.gds1872
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 22.9275 44.466 23.1275 ;
 END
 END vss.gds1872
 PIN vss.gds1873
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 22.9275 43.794 23.1275 ;
 END
 END vss.gds1873
 PIN vss.gds1874
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 22.9275 43.122 23.1275 ;
 END
 END vss.gds1874
 PIN vss.gds1875
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 22.9275 42.45 23.1275 ;
 END
 END vss.gds1875
 PIN vss.gds1876
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 22.9275 41.778 23.1275 ;
 END
 END vss.gds1876
 PIN vss.gds1877
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 22.9275 40.686 23.1275 ;
 END
 END vss.gds1877
 PIN vss.gds1878
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 40.964 24.26 41.02 24.46 ;
 RECT 40.964 23 41.02 23.2 ;
 RECT 40.964 21.74 41.02 21.94 ;
 RECT 40.964 20.48 41.02 20.68 ;
 RECT 40.796 23.07 40.852 23.27 ;
 END
 END vss.gds1878
 PIN vss.gds1879
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 22.122 48.974 22.322 ;
 END
 END vss.gds1879
 PIN vss.gds1880
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 20.862 48.974 21.062 ;
 END
 END vss.gds1880
 PIN vss.gds1881
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 24.642 48.974 24.842 ;
 END
 END vss.gds1881
 PIN vss.gds1882
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 23.382 48.974 23.582 ;
 END
 END vss.gds1882
 PIN vss.gds1883
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 20.822 48.002 21.022 ;
 END
 END vss.gds1883
 PIN vss.gds1884
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 23.342 48.002 23.542 ;
 END
 END vss.gds1884
 PIN vss.gds1885
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 24.602 48.002 24.802 ;
 END
 END vss.gds1885
 PIN vss.gds1886
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 24.84 49.522 25.04 ;
 END
 END vss.gds1886
 PIN vss.gds1887
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.366 24.156 47.422 24.356 ;
 END
 END vss.gds1887
 PIN vss.gds1888
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.254 21.1635 46.314 21.3635 ;
 END
 END vss.gds1888
 PIN vss.gds1889
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.086 21.1635 46.146 21.3635 ;
 END
 END vss.gds1889
 PIN vss.gds1890
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.918 21.1635 45.978 21.3635 ;
 END
 END vss.gds1890
 PIN vss.gds1891
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.582 21.1635 45.642 21.3635 ;
 END
 END vss.gds1891
 PIN vss.gds1892
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.414 21.1635 45.474 21.3635 ;
 END
 END vss.gds1892
 PIN vss.gds1893
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.246 21.1635 45.306 21.3635 ;
 END
 END vss.gds1893
 PIN vss.gds1894
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 22.9275 45.81 23.1275 ;
 END
 END vss.gds1894
 PIN vss.gds1895
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 22.765 46.482 22.965 ;
 END
 END vss.gds1895
 PIN vss.gds1896
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 21.8495 47.162 22.0495 ;
 END
 END vss.gds1896
 PIN vss.gds1897
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 24.097 50.25 24.297 ;
 END
 END vss.gds1897
 PIN vss.gds1898
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 22.837 50.25 23.037 ;
 END
 END vss.gds1898
 PIN vss.gds1899
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 21.577 50.25 21.777 ;
 END
 END vss.gds1899
 PIN vss.gds1900
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 25.357 50.25 25.557 ;
 END
 END vss.gds1900
 PIN vss.gds1901
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 23.0835 46.922 23.2835 ;
 END
 END vss.gds1901
 PIN vss.gds1902
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 23.467 46.694 23.667 ;
 END
 END vss.gds1902
 PIN vss.gds1903
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 22.9275 47.762 23.1275 ;
 END
 END vss.gds1903
 PIN vss.gds1904
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 23.22 49.266 23.42 ;
 END
 END vss.gds1904
 PIN vss.gds1905
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 22.082 48.002 22.282 ;
 END
 END vss.gds1905
 PIN vss.gds1906
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 23.22 48.602 23.42 ;
 END
 END vss.gds1906
 PIN vss.gds1907
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 23.22 49.946 23.42 ;
 END
 END vss.gds1907
 PIN vss.gds1908
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 49.7 21.244 49.756 21.444 ;
 RECT 49.952 21.247 50.008 21.447 ;
 RECT 48.104 22.26 48.16 22.433 ;
 RECT 48.272 22.233 48.328 22.433 ;
 RECT 49.868 22.277 49.924 22.442 ;
 RECT 49.7 22.277 49.756 22.442 ;
 RECT 48.944 22.277 49 22.442 ;
 RECT 48.776 22.277 48.832 22.442 ;
 RECT 48.104 21 48.16 21.173 ;
 RECT 48.272 20.973 48.328 21.173 ;
 RECT 49.868 21.017 49.924 21.182 ;
 RECT 49.7 21.017 49.756 21.182 ;
 RECT 48.944 21.017 49 21.182 ;
 RECT 48.776 21.017 48.832 21.182 ;
 RECT 48.104 23.52 48.16 23.693 ;
 RECT 48.272 23.493 48.328 23.693 ;
 RECT 49.868 23.537 49.924 23.702 ;
 RECT 49.7 23.537 49.756 23.702 ;
 RECT 48.944 23.537 49 23.702 ;
 RECT 48.776 23.537 48.832 23.702 ;
 RECT 49.7 23.764 49.756 23.964 ;
 RECT 49.952 23.767 50.008 23.967 ;
 RECT 48.104 24.78 48.16 24.953 ;
 RECT 48.272 24.753 48.328 24.953 ;
 RECT 49.868 24.797 49.924 24.962 ;
 RECT 49.7 24.797 49.756 24.962 ;
 RECT 48.944 24.797 49 24.962 ;
 RECT 48.776 24.797 48.832 24.962 ;
 RECT 49.7 25.024 49.756 25.224 ;
 RECT 49.952 25.027 50.008 25.227 ;
 RECT 49.7 22.504 49.756 22.704 ;
 RECT 49.952 22.507 50.008 22.707 ;
 RECT 48.44 22.853 48.496 23.053 ;
 RECT 48.272 22.853 48.328 23.053 ;
 RECT 48.44 25.373 48.496 25.573 ;
 RECT 48.272 25.373 48.328 25.573 ;
 RECT 49.112 24.323 49.168 24.523 ;
 RECT 49.532 24.323 49.588 24.523 ;
 RECT 48.44 24.113 48.496 24.313 ;
 RECT 48.272 24.113 48.328 24.313 ;
 RECT 47.768 24.247 47.824 24.447 ;
 RECT 47.768 22.987 47.824 23.187 ;
 RECT 49.112 23.063 49.168 23.263 ;
 RECT 49.532 23.063 49.588 23.263 ;
 RECT 48.44 21.593 48.496 21.793 ;
 RECT 48.272 21.593 48.328 21.793 ;
 RECT 49.112 21.803 49.168 22.003 ;
 RECT 49.532 21.803 49.588 22.003 ;
 RECT 49.112 20.543 49.168 20.743 ;
 RECT 49.532 20.543 49.588 20.743 ;
 RECT 47.768 20.467 47.824 20.667 ;
 RECT 47.768 21.727 47.824 21.927 ;
 RECT 47.6 21.039 47.656 21.239 ;
 RECT 46.928 21.028 46.984 21.228 ;
 RECT 46.592 21.058 46.648 21.258 ;
 RECT 47.432 20.977 47.488 21.177 ;
 RECT 46.76 21.058 46.816 21.258 ;
 RECT 49.28 21.2435 49.336 21.4435 ;
 RECT 47.264 21.028 47.32 21.228 ;
 RECT 47.096 21.028 47.152 21.228 ;
 END
 END vss.gds1908
 PIN vss.gds1909
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.638 21.1635 52.698 21.3635 ;
 END
 END vss.gds1909
 PIN vss.gds1910
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.806 21.1635 52.866 21.3635 ;
 END
 END vss.gds1910
 PIN vss.gds1911
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.142 21.1635 53.202 21.3635 ;
 END
 END vss.gds1911
 PIN vss.gds1912
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.31 21.1635 53.37 21.3635 ;
 END
 END vss.gds1912
 PIN vss.gds1913
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.478 21.1635 53.538 21.3635 ;
 END
 END vss.gds1913
 PIN vss.gds1914
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.814 21.1635 53.874 21.3635 ;
 END
 END vss.gds1914
 PIN vss.gds1915
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.982 21.1635 54.042 21.3635 ;
 END
 END vss.gds1915
 PIN vss.gds1916
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.15 21.1635 54.21 21.3635 ;
 END
 END vss.gds1916
 PIN vss.gds1917
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 22.9275 54.378 23.1275 ;
 END
 END vss.gds1917
 PIN vss.gds1918
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.486 21.1635 54.546 21.3635 ;
 END
 END vss.gds1918
 PIN vss.gds1919
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.654 21.1635 54.714 21.3635 ;
 END
 END vss.gds1919
 PIN vss.gds1920
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.822 21.1635 54.882 21.3635 ;
 END
 END vss.gds1920
 PIN vss.gds1921
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 22.9275 55.05 23.1275 ;
 END
 END vss.gds1921
 PIN vss.gds1922
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.158 21.1635 55.218 21.3635 ;
 END
 END vss.gds1922
 PIN vss.gds1923
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 21.636 50.918 21.836 ;
 END
 END vss.gds1923
 PIN vss.gds1924
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.542 23.7395 51.598 23.9395 ;
 END
 END vss.gds1924
 PIN vss.gds1925
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 22.9275 53.706 23.1275 ;
 END
 END vss.gds1925
 PIN vss.gds1926
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.47 21.1635 52.53 21.3635 ;
 END
 END vss.gds1926
 PIN vss.gds1927
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 24.8475 51.418 25.0475 ;
 END
 END vss.gds1927
 PIN vss.gds1928
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 22.9275 53.034 23.1275 ;
 END
 END vss.gds1928
 PIN vss.gds1929
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.09 20.947 52.13 21.147 ;
 END
 END vss.gds1929
 PIN vss.gds1930
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 23.0835 51.938 23.2835 ;
 END
 END vss.gds1930
 PIN vss.gds1931
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 23.4905 50.594 23.6905 ;
 END
 END vss.gds1931
 PIN vss.gds1932
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 22.765 52.362 22.965 ;
 END
 END vss.gds1932
 PIN vss.gds1933
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 22.8865 51.098 23.0865 ;
 END
 END vss.gds1933
 PIN vss.gds1934
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 50.624 22.28 50.68 22.433 ;
 RECT 50.624 21.02 50.68 21.173 ;
 RECT 50.624 23.54 50.68 23.693 ;
 RECT 50.624 24.8 50.68 24.953 ;
 RECT 50.96 25.4315 51.016 25.6315 ;
 RECT 50.96 24.1715 51.016 24.3715 ;
 RECT 50.456 24.4235 50.512 24.6235 ;
 RECT 50.456 23.1635 50.512 23.3635 ;
 RECT 50.96 22.9115 51.016 23.1115 ;
 RECT 50.456 21.9035 50.512 22.1035 ;
 RECT 50.96 21.6515 51.016 21.8515 ;
 RECT 50.456 20.6435 50.512 20.8435 ;
 RECT 51.968 21.058 52.024 21.258 ;
 RECT 51.8 21.0655 51.856 21.2655 ;
 RECT 51.632 21.058 51.688 21.258 ;
 RECT 51.464 21.058 51.52 21.258 ;
 RECT 51.296 21.058 51.352 21.258 ;
 RECT 51.128 21.173 51.184 21.373 ;
 RECT 52.136 21.058 52.192 21.258 ;
 END
 END vss.gds1934
 PIN vss.gds1935
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 22.9275 60.174 23.1275 ;
 END
 END vss.gds1935
 PIN vss.gds1936
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.946 21.1635 60.006 21.3635 ;
 END
 END vss.gds1936
 PIN vss.gds1937
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.778 21.1635 59.838 21.3635 ;
 END
 END vss.gds1937
 PIN vss.gds1938
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.61 21.1635 59.67 21.3635 ;
 END
 END vss.gds1938
 PIN vss.gds1939
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 22.9275 59.502 23.1275 ;
 END
 END vss.gds1939
 PIN vss.gds1940
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.274 21.1635 59.334 21.3635 ;
 END
 END vss.gds1940
 PIN vss.gds1941
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.106 21.1635 59.166 21.3635 ;
 END
 END vss.gds1941
 PIN vss.gds1942
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.938 21.1635 58.998 21.3635 ;
 END
 END vss.gds1942
 PIN vss.gds1943
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 22.9275 58.83 23.1275 ;
 END
 END vss.gds1943
 PIN vss.gds1944
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.602 21.1635 58.662 21.3635 ;
 END
 END vss.gds1944
 PIN vss.gds1945
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.434 21.1635 58.494 21.3635 ;
 END
 END vss.gds1945
 PIN vss.gds1946
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.266 21.1635 58.326 21.3635 ;
 END
 END vss.gds1946
 PIN vss.gds1947
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.326 21.1635 55.386 21.3635 ;
 END
 END vss.gds1947
 PIN vss.gds1948
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.494 21.1635 55.554 21.3635 ;
 END
 END vss.gds1948
 PIN vss.gds1949
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 22.9275 55.722 23.1275 ;
 END
 END vss.gds1949
 PIN vss.gds1950
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.83 21.1635 55.89 21.3635 ;
 END
 END vss.gds1950
 PIN vss.gds1951
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.998 21.1635 56.058 21.3635 ;
 END
 END vss.gds1951
 PIN vss.gds1952
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.166 21.1635 56.226 21.3635 ;
 END
 END vss.gds1952
 PIN vss.gds1953
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.502 21.1635 56.562 21.3635 ;
 END
 END vss.gds1953
 PIN vss.gds1954
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.67 21.1635 56.73 21.3635 ;
 END
 END vss.gds1954
 PIN vss.gds1955
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.838 21.1635 56.898 21.3635 ;
 END
 END vss.gds1955
 PIN vss.gds1956
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.342 21.1635 57.402 21.3635 ;
 END
 END vss.gds1956
 PIN vss.gds1957
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.51 21.1635 57.57 21.3635 ;
 END
 END vss.gds1957
 PIN vss.gds1958
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.174 21.1635 57.234 21.3635 ;
 END
 END vss.gds1958
 PIN vss.gds1959
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 22.9275 56.394 23.1275 ;
 END
 END vss.gds1959
 PIN vss.gds1960
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 22.9275 57.738 23.1275 ;
 END
 END vss.gds1960
 PIN vss.gds1961
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 22.9275 57.066 23.1275 ;
 END
 END vss.gds1961
 PIN vss.gds1962
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 58.016 23 58.072 23.2 ;
 RECT 58.016 24.26 58.072 24.46 ;
 RECT 58.016 21.74 58.072 21.94 ;
 RECT 58.016 20.48 58.072 20.68 ;
 RECT 57.848 23.07 57.904 23.27 ;
 END
 END vss.gds1962
 PIN vss.gds1963
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 20.822 65.054 21.022 ;
 END
 END vss.gds1963
 PIN vss.gds1964
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 23.342 65.054 23.542 ;
 END
 END vss.gds1964
 PIN vss.gds1965
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 24.602 65.054 24.802 ;
 END
 END vss.gds1965
 PIN vss.gds1966
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 21.8495 64.214 22.0495 ;
 END
 END vss.gds1966
 PIN vss.gds1967
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.418 24.156 64.474 24.356 ;
 END
 END vss.gds1967
 PIN vss.gds1968
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 22.765 63.534 22.965 ;
 END
 END vss.gds1968
 PIN vss.gds1969
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.306 21.1635 63.366 21.3635 ;
 END
 END vss.gds1969
 PIN vss.gds1970
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.138 21.1635 63.198 21.3635 ;
 END
 END vss.gds1970
 PIN vss.gds1971
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.97 21.1635 63.03 21.3635 ;
 END
 END vss.gds1971
 PIN vss.gds1972
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 22.9275 62.862 23.1275 ;
 END
 END vss.gds1972
 PIN vss.gds1973
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.634 21.1635 62.694 21.3635 ;
 END
 END vss.gds1973
 PIN vss.gds1974
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.466 21.1635 62.526 21.3635 ;
 END
 END vss.gds1974
 PIN vss.gds1975
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.298 21.1635 62.358 21.3635 ;
 END
 END vss.gds1975
 PIN vss.gds1976
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 22.9275 62.19 23.1275 ;
 END
 END vss.gds1976
 PIN vss.gds1977
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.962 21.1635 62.022 21.3635 ;
 END
 END vss.gds1977
 PIN vss.gds1978
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.794 21.1635 61.854 21.3635 ;
 END
 END vss.gds1978
 PIN vss.gds1979
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.626 21.1635 61.686 21.3635 ;
 END
 END vss.gds1979
 PIN vss.gds1980
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 22.9275 61.518 23.1275 ;
 END
 END vss.gds1980
 PIN vss.gds1981
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.29 21.1635 61.35 21.3635 ;
 END
 END vss.gds1981
 PIN vss.gds1982
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.122 21.1635 61.182 21.3635 ;
 END
 END vss.gds1982
 PIN vss.gds1983
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.954 21.1635 61.014 21.3635 ;
 END
 END vss.gds1983
 PIN vss.gds1984
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 22.9275 60.846 23.1275 ;
 END
 END vss.gds1984
 PIN vss.gds1985
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.618 21.1635 60.678 21.3635 ;
 END
 END vss.gds1985
 PIN vss.gds1986
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.45 21.1635 60.51 21.3635 ;
 END
 END vss.gds1986
 PIN vss.gds1987
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.282 21.1635 60.342 21.3635 ;
 END
 END vss.gds1987
 PIN vss.gds1988
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 22.082 65.054 22.282 ;
 END
 END vss.gds1988
 PIN vss.gds1989
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 23.0835 63.974 23.2835 ;
 END
 END vss.gds1989
 PIN vss.gds1990
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 23.467 63.746 23.667 ;
 END
 END vss.gds1990
 PIN vss.gds1991
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 22.9275 64.814 23.1275 ;
 END
 END vss.gds1991
 PIN vss.gds1992
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 65.156 22.26 65.212 22.433 ;
 RECT 65.156 21 65.212 21.173 ;
 RECT 65.156 23.52 65.212 23.693 ;
 RECT 65.156 24.78 65.212 24.953 ;
 RECT 64.82 24.247 64.876 24.447 ;
 RECT 64.82 22.987 64.876 23.187 ;
 RECT 64.82 21.727 64.876 21.927 ;
 RECT 64.82 20.467 64.876 20.667 ;
 RECT 64.652 21.039 64.708 21.239 ;
 RECT 63.98 21.028 64.036 21.228 ;
 RECT 64.484 20.977 64.54 21.177 ;
 RECT 63.812 21.058 63.868 21.258 ;
 RECT 64.316 21.028 64.372 21.228 ;
 RECT 64.148 21.028 64.204 21.228 ;
 RECT 63.644 21.058 63.7 21.258 ;
 END
 END vss.gds1992
 PIN vss.gds1993
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 22.122 66.026 22.322 ;
 END
 END vss.gds1993
 PIN vss.gds1994
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 20.862 66.026 21.062 ;
 END
 END vss.gds1994
 PIN vss.gds1995
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 24.642 66.026 24.842 ;
 END
 END vss.gds1995
 PIN vss.gds1996
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 23.382 66.026 23.582 ;
 END
 END vss.gds1996
 PIN vss.gds1997
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 24.097 67.302 24.297 ;
 END
 END vss.gds1997
 PIN vss.gds1998
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 23.22 66.318 23.42 ;
 END
 END vss.gds1998
 PIN vss.gds1999
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 24.84 66.574 25.04 ;
 END
 END vss.gds1999
 PIN vss.gds2000
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.142 20.947 69.182 21.147 ;
 END
 END vss.gds2000
 PIN vss.gds2001
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.69 21.1635 69.75 21.3635 ;
 END
 END vss.gds2001
 PIN vss.gds2002
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.858 21.1635 69.918 21.3635 ;
 END
 END vss.gds2002
 PIN vss.gds2003
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 22.9275 70.086 23.1275 ;
 END
 END vss.gds2003
 PIN vss.gds2004
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.194 21.1635 70.254 21.3635 ;
 END
 END vss.gds2004
 PIN vss.gds2005
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.594 23.7395 68.65 23.9395 ;
 END
 END vss.gds2005
 PIN vss.gds2006
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 21.636 67.97 21.836 ;
 END
 END vss.gds2006
 PIN vss.gds2007
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 25.357 67.302 25.557 ;
 END
 END vss.gds2007
 PIN vss.gds2008
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 22.837 67.302 23.037 ;
 END
 END vss.gds2008
 PIN vss.gds2009
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 21.577 67.302 21.777 ;
 END
 END vss.gds2009
 PIN vss.gds2010
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.522 21.1635 69.582 21.3635 ;
 END
 END vss.gds2010
 PIN vss.gds2011
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 22.8865 68.15 23.0865 ;
 END
 END vss.gds2011
 PIN vss.gds2012
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 24.8475 68.47 25.0475 ;
 END
 END vss.gds2012
 PIN vss.gds2013
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 23.4905 67.646 23.6905 ;
 END
 END vss.gds2013
 PIN vss.gds2014
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 23.22 65.654 23.42 ;
 END
 END vss.gds2014
 PIN vss.gds2015
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 23.22 66.998 23.42 ;
 END
 END vss.gds2015
 PIN vss.gds2016
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 23.0835 68.99 23.2835 ;
 END
 END vss.gds2016
 PIN vss.gds2017
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 22.765 69.414 22.965 ;
 END
 END vss.gds2017
 PIN vss.gds2018
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 66.752 21.244 66.808 21.444 ;
 RECT 67.004 21.247 67.06 21.447 ;
 RECT 67.676 22.28 67.732 22.433 ;
 RECT 65.324 22.233 65.38 22.433 ;
 RECT 66.92 22.277 66.976 22.442 ;
 RECT 66.752 22.277 66.808 22.442 ;
 RECT 65.996 22.277 66.052 22.442 ;
 RECT 65.828 22.277 65.884 22.442 ;
 RECT 67.676 21.02 67.732 21.173 ;
 RECT 65.324 20.973 65.38 21.173 ;
 RECT 66.92 21.017 66.976 21.182 ;
 RECT 66.752 21.017 66.808 21.182 ;
 RECT 65.996 21.017 66.052 21.182 ;
 RECT 65.828 21.017 65.884 21.182 ;
 RECT 67.676 23.54 67.732 23.693 ;
 RECT 65.324 23.493 65.38 23.693 ;
 RECT 66.92 23.537 66.976 23.702 ;
 RECT 66.752 23.537 66.808 23.702 ;
 RECT 65.996 23.537 66.052 23.702 ;
 RECT 65.828 23.537 65.884 23.702 ;
 RECT 67.676 24.8 67.732 24.953 ;
 RECT 65.324 24.753 65.38 24.953 ;
 RECT 66.92 24.797 66.976 24.962 ;
 RECT 66.752 24.797 66.808 24.962 ;
 RECT 65.996 24.797 66.052 24.962 ;
 RECT 65.828 24.797 65.884 24.962 ;
 RECT 66.752 22.504 66.808 22.704 ;
 RECT 67.004 22.507 67.06 22.707 ;
 RECT 66.752 23.764 66.808 23.964 ;
 RECT 67.004 23.767 67.06 23.967 ;
 RECT 66.752 25.024 66.808 25.224 ;
 RECT 67.004 25.027 67.06 25.227 ;
 RECT 66.164 24.323 66.22 24.523 ;
 RECT 65.492 24.113 65.548 24.313 ;
 RECT 65.324 24.113 65.38 24.313 ;
 RECT 68.012 24.1715 68.068 24.3715 ;
 RECT 67.508 24.4235 67.564 24.6235 ;
 RECT 68.012 25.4315 68.068 25.6315 ;
 RECT 65.492 25.373 65.548 25.573 ;
 RECT 65.324 25.373 65.38 25.573 ;
 RECT 66.584 24.323 66.64 24.523 ;
 RECT 65.492 21.593 65.548 21.793 ;
 RECT 65.324 21.593 65.38 21.793 ;
 RECT 66.164 21.803 66.22 22.003 ;
 RECT 66.584 21.803 66.64 22.003 ;
 RECT 68.012 22.9115 68.068 23.1115 ;
 RECT 67.508 23.1635 67.564 23.3635 ;
 RECT 66.164 23.063 66.22 23.263 ;
 RECT 66.584 23.063 66.64 23.263 ;
 RECT 65.492 22.853 65.548 23.053 ;
 RECT 65.324 22.853 65.38 23.053 ;
 RECT 67.508 21.9035 67.564 22.1035 ;
 RECT 68.012 21.6515 68.068 21.8515 ;
 RECT 66.164 20.543 66.22 20.743 ;
 RECT 66.584 20.543 66.64 20.743 ;
 RECT 67.508 20.6435 67.564 20.8435 ;
 RECT 66.332 21.2435 66.388 21.4435 ;
 RECT 69.02 21.058 69.076 21.258 ;
 RECT 68.852 21.0655 68.908 21.2655 ;
 RECT 68.684 21.058 68.74 21.258 ;
 RECT 68.516 21.058 68.572 21.258 ;
 RECT 68.348 21.058 68.404 21.258 ;
 RECT 69.188 21.058 69.244 21.258 ;
 RECT 68.18 21.173 68.236 21.373 ;
 END
 END vss.gds2018
 PIN vss.gds2019
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.362 21.1635 70.422 21.3635 ;
 END
 END vss.gds2019
 PIN vss.gds2020
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.53 21.1635 70.59 21.3635 ;
 END
 END vss.gds2020
 PIN vss.gds2021
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.866 21.1635 70.926 21.3635 ;
 END
 END vss.gds2021
 PIN vss.gds2022
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.034 21.1635 71.094 21.3635 ;
 END
 END vss.gds2022
 PIN vss.gds2023
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.202 21.1635 71.262 21.3635 ;
 END
 END vss.gds2023
 PIN vss.gds2024
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 22.9275 71.43 23.1275 ;
 END
 END vss.gds2024
 PIN vss.gds2025
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.538 21.1635 71.598 21.3635 ;
 END
 END vss.gds2025
 PIN vss.gds2026
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.706 21.1635 71.766 21.3635 ;
 END
 END vss.gds2026
 PIN vss.gds2027
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.874 21.1635 71.934 21.3635 ;
 END
 END vss.gds2027
 PIN vss.gds2028
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 22.9275 72.102 23.1275 ;
 END
 END vss.gds2028
 PIN vss.gds2029
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.21 21.1635 72.27 21.3635 ;
 END
 END vss.gds2029
 PIN vss.gds2030
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.378 21.1635 72.438 21.3635 ;
 END
 END vss.gds2030
 PIN vss.gds2031
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.546 21.1635 72.606 21.3635 ;
 END
 END vss.gds2031
 PIN vss.gds2032
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 22.9275 72.774 23.1275 ;
 END
 END vss.gds2032
 PIN vss.gds2033
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.882 21.1635 72.942 21.3635 ;
 END
 END vss.gds2033
 PIN vss.gds2034
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.05 21.1635 73.11 21.3635 ;
 END
 END vss.gds2034
 PIN vss.gds2035
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.554 21.1635 73.614 21.3635 ;
 END
 END vss.gds2035
 PIN vss.gds2036
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.722 21.1635 73.782 21.3635 ;
 END
 END vss.gds2036
 PIN vss.gds2037
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.89 21.1635 73.95 21.3635 ;
 END
 END vss.gds2037
 PIN vss.gds2038
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.226 21.1635 74.286 21.3635 ;
 END
 END vss.gds2038
 PIN vss.gds2039
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.394 21.1635 74.454 21.3635 ;
 END
 END vss.gds2039
 PIN vss.gds2040
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.218 21.1635 73.278 21.3635 ;
 END
 END vss.gds2040
 PIN vss.gds2041
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.562 21.1635 74.622 21.3635 ;
 END
 END vss.gds2041
 PIN vss.gds2042
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 22.9275 70.758 23.1275 ;
 END
 END vss.gds2042
 PIN vss.gds2043
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 22.9275 74.118 23.1275 ;
 END
 END vss.gds2043
 PIN vss.gds2044
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 22.9275 74.79 23.1275 ;
 END
 END vss.gds2044
 PIN vss.gds2045
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 22.9275 73.446 23.1275 ;
 END
 END vss.gds2045
 PIN vss.gds2046
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 27.7925 0.29 27.9925 ;
 END
 END vss.gds2046
 PIN vss.gds2047
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 27.877 2.962 28.077 ;
 END
 END vss.gds2047
 PIN vss.gds2048
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 26.617 2.962 26.817 ;
 END
 END vss.gds2048
 PIN vss.gds2049
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.286 25.987 3.326 26.187 ;
 END
 END vss.gds2049
 PIN vss.gds2050
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 27.476 3.142 27.676 ;
 END
 END vss.gds2050
 PIN vss.gds2051
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 26.216 3.142 26.416 ;
 END
 END vss.gds2051
 PIN vss.gds2052
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.442 25.581 4.482 25.781 ;
 END
 END vss.gds2052
 PIN vss.gds2053
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.414 26.263 3.454 26.463 ;
 END
 END vss.gds2053
 PIN vss.gds2054
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 27.042 0.602 27.242 ;
 END
 END vss.gds2054
 PIN vss.gds2055
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 26.841 0.942 27.041 ;
 END
 END vss.gds2055
 PIN vss.gds2056
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 27.385 1.282 27.585 ;
 END
 END vss.gds2056
 PIN vss.gds2057
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 27.2705 2.122 27.4705 ;
 END
 END vss.gds2057
 PIN vss.gds2058
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.754 27.247 3.794 27.447 ;
 END
 END vss.gds2058
 PIN vss.gds2059
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 27.247 5.074 27.447 ;
 END
 END vss.gds2059
 PIN vss.gds2060
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 27.247 4.194 27.447 ;
 END
 END vss.gds2060
 PIN vss.gds2061
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 28.566 3.142 28.766 ;
 END
 END vss.gds2061
 PIN vss.gds2062
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.57 25.784 4.61 25.984 ;
 END
 END vss.gds2062
 PIN vss.gds2063
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 25.581 4.882 25.781 ;
 END
 END vss.gds2063
 PIN vss.gds2064
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 27.1435 4.002 27.3435 ;
 END
 END vss.gds2064
 PIN vss.gds2065
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 27.1435 5.282 27.3435 ;
 END
 END vss.gds2065
 PIN vss.gds2066
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.562 26.263 3.602 26.463 ;
 END
 END vss.gds2066
 PIN vss.gds2067
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 26.872 2.302 27.072 ;
 END
 END vss.gds2067
 PIN vss.gds2068
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 27.442 1.462 27.642 ;
 END
 END vss.gds2068
 PIN vss.gds2069
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 26.9415 0.718 27.1415 ;
 END
 END vss.gds2069
 PIN vss.gds2070
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 3.332 25.449 3.388 25.649 ;
 RECT 2.576 26.6175 2.632 26.8175 ;
 RECT 2.408 26.6175 2.464 26.8175 ;
 RECT 2.996 26.6175 3.052 26.8175 ;
 RECT 3.332 26.709 3.388 26.909 ;
 RECT 3.5 26.6655 3.556 26.8655 ;
 RECT 0.98 26.5325 1.036 26.7325 ;
 RECT 2.072 26.533 2.128 26.733 ;
 RECT 2.576 27.8775 2.632 28.0775 ;
 RECT 2.408 27.8775 2.464 28.0775 ;
 RECT 2.996 27.8775 3.052 28.0775 ;
 RECT 3.332 27.969 3.388 28.169 ;
 RECT 3.5 27.9255 3.556 28.1255 ;
 RECT 0.98 27.7925 1.036 27.9925 ;
 RECT 2.072 27.793 2.128 27.993 ;
 RECT 0.392 27.883 0.448 28.083 ;
 RECT 0.812 27.969 0.868 28.169 ;
 RECT 0.644 27.883 0.7 28.083 ;
 RECT 1.232 27.883 1.288 28.083 ;
 RECT 1.4 27.883 1.456 28.083 ;
 RECT 1.568 27.883 1.624 28.083 ;
 RECT 1.82 27.883 1.876 28.083 ;
 RECT 2.24 27.883 2.296 28.083 ;
 RECT 2.744 27.793 2.8 27.993 ;
 RECT 3.164 27.883 3.22 28.083 ;
 RECT 3.92 27.883 3.976 28.083 ;
 RECT 3.752 28.153 3.808 28.353 ;
 RECT 4.508 28.0825 4.564 28.2825 ;
 RECT 0.392 26.623 0.448 26.823 ;
 RECT 0.812 26.709 0.868 26.909 ;
 RECT 0.644 26.623 0.7 26.823 ;
 RECT 1.232 26.623 1.288 26.823 ;
 RECT 1.4 26.623 1.456 26.823 ;
 RECT 1.568 26.623 1.624 26.823 ;
 RECT 1.82 26.623 1.876 26.823 ;
 RECT 2.24 26.623 2.296 26.823 ;
 RECT 2.744 26.533 2.8 26.733 ;
 RECT 3.164 26.623 3.22 26.823 ;
 RECT 3.92 26.623 3.976 26.823 ;
 RECT 3.752 26.893 3.808 27.093 ;
 RECT 4.508 26.8225 4.564 27.0225 ;
 RECT 0.812 25.449 0.868 25.649 ;
 RECT 3.752 25.633 3.808 25.833 ;
 RECT 4.508 25.5625 4.564 25.7625 ;
 END
 END vss.gds2070
 PIN vss.gds2071
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.134 26.2035 10.194 26.4035 ;
 END
 END vss.gds2071
 PIN vss.gds2072
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.966 26.2035 10.026 26.4035 ;
 END
 END vss.gds2072
 PIN vss.gds2073
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.798 26.2035 9.858 26.4035 ;
 END
 END vss.gds2073
 PIN vss.gds2074
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.462 26.2035 9.522 26.4035 ;
 END
 END vss.gds2074
 PIN vss.gds2075
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.294 26.2035 9.354 26.4035 ;
 END
 END vss.gds2075
 PIN vss.gds2076
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.79 26.2035 8.85 26.4035 ;
 END
 END vss.gds2076
 PIN vss.gds2077
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.622 26.2035 8.682 26.4035 ;
 END
 END vss.gds2077
 PIN vss.gds2078
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.454 26.2035 8.514 26.4035 ;
 END
 END vss.gds2078
 PIN vss.gds2079
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.118 26.2035 8.178 26.4035 ;
 END
 END vss.gds2079
 PIN vss.gds2080
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.95 26.2035 8.01 26.4035 ;
 END
 END vss.gds2080
 PIN vss.gds2081
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.782 26.2035 7.842 26.4035 ;
 END
 END vss.gds2081
 PIN vss.gds2082
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.126 26.2035 9.186 26.4035 ;
 END
 END vss.gds2082
 PIN vss.gds2083
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.446 26.2035 7.506 26.4035 ;
 END
 END vss.gds2083
 PIN vss.gds2084
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.278 26.2035 7.338 26.4035 ;
 END
 END vss.gds2084
 PIN vss.gds2085
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 27.092 9.69 27.292 ;
 END
 END vss.gds2085
 PIN vss.gds2086
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 27.092 8.346 27.292 ;
 END
 END vss.gds2086
 PIN vss.gds2087
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 27.092 9.018 27.292 ;
 END
 END vss.gds2087
 PIN vss.gds2088
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 27.092 7.674 27.292 ;
 END
 END vss.gds2088
 PIN vss.gds2089
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.11 26.2035 7.17 26.4035 ;
 END
 END vss.gds2089
 PIN vss.gds2090
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 27.247 5.474 27.447 ;
 END
 END vss.gds2090
 PIN vss.gds2091
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 27.247 5.986 27.447 ;
 END
 END vss.gds2091
 PIN vss.gds2092
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 27.044 6.178 27.244 ;
 END
 END vss.gds2092
 PIN vss.gds2093
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 27.247 5.73 27.447 ;
 END
 END vss.gds2093
 PIN vss.gds2094
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 27.043 6.434 27.243 ;
 END
 END vss.gds2094
 PIN vss.gds2095
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 6.524 26.585 6.58 26.785 ;
 RECT 6.524 27.845 6.58 28.045 ;
 RECT 6.692 25.648 6.748 25.848 ;
 RECT 6.692 26.908 6.748 27.108 ;
 RECT 6.692 28.168 6.748 28.368 ;
 RECT 6.608 28.153 6.664 28.353 ;
 RECT 6.608 26.893 6.664 27.093 ;
 RECT 6.608 25.633 6.664 25.833 ;
 END
 END vss.gds2095
 PIN vss.gds2096
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 28.382 13.898 28.582 ;
 END
 END vss.gds2096
 PIN vss.gds2097
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 28.422 14.87 28.622 ;
 END
 END vss.gds2097
 PIN vss.gds2098
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 25.862 13.898 26.062 ;
 END
 END vss.gds2098
 PIN vss.gds2099
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 25.902 14.87 26.102 ;
 END
 END vss.gds2099
 PIN vss.gds2100
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 27.122 13.898 27.322 ;
 END
 END vss.gds2100
 PIN vss.gds2101
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 27.162 14.87 27.362 ;
 END
 END vss.gds2101
 PIN vss.gds2102
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.15 26.2035 12.21 26.4035 ;
 END
 END vss.gds2102
 PIN vss.gds2103
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.982 26.2035 12.042 26.4035 ;
 END
 END vss.gds2103
 PIN vss.gds2104
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.814 26.2035 11.874 26.4035 ;
 END
 END vss.gds2104
 PIN vss.gds2105
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.478 26.2035 11.538 26.4035 ;
 END
 END vss.gds2105
 PIN vss.gds2106
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.31 26.2035 11.37 26.4035 ;
 END
 END vss.gds2106
 PIN vss.gds2107
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.142 26.2035 11.202 26.4035 ;
 END
 END vss.gds2107
 PIN vss.gds2108
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.806 26.2035 10.866 26.4035 ;
 END
 END vss.gds2108
 PIN vss.gds2109
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.638 26.2035 10.698 26.4035 ;
 END
 END vss.gds2109
 PIN vss.gds2110
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.47 26.2035 10.53 26.4035 ;
 END
 END vss.gds2110
 PIN vss.gds2111
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 27.092 13.658 27.292 ;
 END
 END vss.gds2111
 PIN vss.gds2112
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 26.568 13.058 26.768 ;
 END
 END vss.gds2112
 PIN vss.gds2113
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.262 27.777 13.318 27.977 ;
 END
 END vss.gds2113
 PIN vss.gds2114
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 27.092 11.706 27.292 ;
 END
 END vss.gds2114
 PIN vss.gds2115
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 27.092 11.034 27.292 ;
 END
 END vss.gds2115
 PIN vss.gds2116
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 27.247 15.162 27.447 ;
 END
 END vss.gds2116
 PIN vss.gds2117
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 27.092 10.362 27.292 ;
 END
 END vss.gds2117
 PIN vss.gds2118
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 27.247 14.498 27.447 ;
 END
 END vss.gds2118
 PIN vss.gds2119
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 27.1335 12.818 27.3335 ;
 END
 END vss.gds2119
 PIN vss.gds2120
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 26.9805 12.378 27.1805 ;
 END
 END vss.gds2120
 PIN vss.gds2121
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 27.247 12.59 27.447 ;
 END
 END vss.gds2121
 PIN vss.gds2122
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 14 28.56 14.056 28.733 ;
 RECT 14.168 28.533 14.224 28.733 ;
 RECT 14 27.3 14.056 27.473 ;
 RECT 14.168 27.273 14.224 27.473 ;
 RECT 14 26.04 14.056 26.213 ;
 RECT 14.168 26.013 14.224 26.213 ;
 RECT 14.336 26.633 14.392 26.833 ;
 RECT 14.168 26.633 14.224 26.833 ;
 RECT 15.008 25.583 15.064 25.783 ;
 RECT 14.84 26.057 14.896 26.222 ;
 RECT 14.672 26.057 14.728 26.222 ;
 RECT 13.664 25.507 13.72 25.707 ;
 RECT 15.008 26.843 15.064 27.043 ;
 RECT 14.84 27.317 14.896 27.482 ;
 RECT 14.672 27.317 14.728 27.482 ;
 RECT 13.664 26.767 13.72 26.967 ;
 RECT 15.008 28.103 15.064 28.303 ;
 RECT 14.84 28.577 14.896 28.742 ;
 RECT 14.672 28.577 14.728 28.742 ;
 RECT 14.336 27.893 14.392 28.093 ;
 RECT 14.168 27.893 14.224 28.093 ;
 RECT 13.664 28.027 13.72 28.227 ;
 RECT 15.176 26.2835 15.232 26.4835 ;
 RECT 12.824 28.67 12.88 28.87 ;
 RECT 12.824 26.068 12.88 26.268 ;
 RECT 13.496 26.079 13.552 26.279 ;
 RECT 13.328 28.67 13.384 28.87 ;
 RECT 13.328 26.017 13.384 26.217 ;
 RECT 13.16 28.67 13.216 28.87 ;
 RECT 13.16 26.068 13.216 26.268 ;
 RECT 12.488 28.67 12.544 28.87 ;
 RECT 12.488 26.098 12.544 26.298 ;
 RECT 12.992 28.67 13.048 28.87 ;
 RECT 12.992 26.068 13.048 26.268 ;
 RECT 12.656 28.67 12.712 28.87 ;
 RECT 12.656 26.098 12.712 26.298 ;
 END
 END vss.gds2122
 PIN vss.gds2123
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.986 25.987 18.026 26.187 ;
 END
 END vss.gds2123
 PIN vss.gds2124
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 27.99 15.418 28.19 ;
 END
 END vss.gds2124
 PIN vss.gds2125
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.438 27.5195 17.494 27.7195 ;
 END
 END vss.gds2125
 PIN vss.gds2126
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.038 26.2035 19.098 26.4035 ;
 END
 END vss.gds2126
 PIN vss.gds2127
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.206 26.2035 19.266 26.4035 ;
 END
 END vss.gds2127
 PIN vss.gds2128
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.374 26.2035 19.434 26.4035 ;
 END
 END vss.gds2128
 PIN vss.gds2129
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 27.092 20.274 27.292 ;
 END
 END vss.gds2129
 PIN vss.gds2130
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 27.877 16.146 28.077 ;
 END
 END vss.gds2130
 PIN vss.gds2131
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 26.617 16.146 26.817 ;
 END
 END vss.gds2131
 PIN vss.gds2132
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.702 26.2035 18.762 26.4035 ;
 END
 END vss.gds2132
 PIN vss.gds2133
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.71 26.2035 19.77 26.4035 ;
 END
 END vss.gds2133
 PIN vss.gds2134
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.878 26.2035 19.938 26.4035 ;
 END
 END vss.gds2134
 PIN vss.gds2135
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.534 26.2035 18.594 26.4035 ;
 END
 END vss.gds2135
 PIN vss.gds2136
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 26.4895 16.814 26.6895 ;
 END
 END vss.gds2136
 PIN vss.gds2137
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 27.9975 17.314 28.1975 ;
 END
 END vss.gds2137
 PIN vss.gds2138
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.366 26.2035 18.426 26.4035 ;
 END
 END vss.gds2138
 PIN vss.gds2139
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.046 26.2035 20.106 26.4035 ;
 END
 END vss.gds2139
 PIN vss.gds2140
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 27.092 19.602 27.292 ;
 END
 END vss.gds2140
 PIN vss.gds2141
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 27.092 18.93 27.292 ;
 END
 END vss.gds2141
 PIN vss.gds2142
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 27.0605 16.994 27.2605 ;
 END
 END vss.gds2142
 PIN vss.gds2143
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 27.247 15.842 27.447 ;
 END
 END vss.gds2143
 PIN vss.gds2144
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 27.1335 17.834 27.3335 ;
 END
 END vss.gds2144
 PIN vss.gds2145
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 27.2705 16.49 27.4705 ;
 END
 END vss.gds2145
 PIN vss.gds2146
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 26.9805 18.258 27.1805 ;
 END
 END vss.gds2146
 PIN vss.gds2147
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 15.596 27.544 15.652 27.744 ;
 RECT 15.848 27.547 15.904 27.747 ;
 RECT 16.52 28.58 16.576 28.733 ;
 RECT 15.764 28.577 15.82 28.742 ;
 RECT 15.596 28.577 15.652 28.742 ;
 RECT 15.596 26.284 15.652 26.484 ;
 RECT 15.848 26.287 15.904 26.487 ;
 RECT 16.52 27.32 16.576 27.473 ;
 RECT 15.764 27.317 15.82 27.482 ;
 RECT 15.596 27.317 15.652 27.482 ;
 RECT 16.52 26.06 16.576 26.213 ;
 RECT 15.764 26.057 15.82 26.222 ;
 RECT 15.596 26.057 15.652 26.222 ;
 RECT 15.428 25.583 15.484 25.783 ;
 RECT 16.352 25.6835 16.408 25.8835 ;
 RECT 15.428 26.843 15.484 27.043 ;
 RECT 16.352 26.9435 16.408 27.1435 ;
 RECT 16.856 26.6915 16.912 26.8915 ;
 RECT 16.856 27.9515 16.912 28.1515 ;
 RECT 16.352 28.2035 16.408 28.4035 ;
 RECT 15.428 28.103 15.484 28.303 ;
 RECT 17.864 28.67 17.92 28.87 ;
 RECT 17.864 26.098 17.92 26.298 ;
 RECT 17.696 28.67 17.752 28.87 ;
 RECT 17.696 26.1055 17.752 26.3055 ;
 RECT 17.528 28.67 17.584 28.87 ;
 RECT 17.528 26.098 17.584 26.298 ;
 RECT 17.36 28.67 17.416 28.87 ;
 RECT 17.36 26.098 17.416 26.298 ;
 RECT 17.192 28.67 17.248 28.87 ;
 RECT 17.192 26.098 17.248 26.298 ;
 RECT 18.032 28.67 18.088 28.87 ;
 RECT 18.032 26.098 18.088 26.298 ;
 RECT 17.024 26.213 17.08 26.413 ;
 END
 END vss.gds2147
 PIN vss.gds2148
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.17 26.2035 25.23 26.4035 ;
 END
 END vss.gds2148
 PIN vss.gds2149
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.002 26.2035 25.062 26.4035 ;
 END
 END vss.gds2149
 PIN vss.gds2150
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.834 26.2035 24.894 26.4035 ;
 END
 END vss.gds2150
 PIN vss.gds2151
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.498 26.2035 24.558 26.4035 ;
 END
 END vss.gds2151
 PIN vss.gds2152
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.33 26.2035 24.39 26.4035 ;
 END
 END vss.gds2152
 PIN vss.gds2153
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.162 26.2035 24.222 26.4035 ;
 END
 END vss.gds2153
 PIN vss.gds2154
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.382 26.2035 20.442 26.4035 ;
 END
 END vss.gds2154
 PIN vss.gds2155
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.55 26.2035 20.61 26.4035 ;
 END
 END vss.gds2155
 PIN vss.gds2156
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.718 26.2035 20.778 26.4035 ;
 END
 END vss.gds2156
 PIN vss.gds2157
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.054 26.2035 21.114 26.4035 ;
 END
 END vss.gds2157
 PIN vss.gds2158
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.222 26.2035 21.282 26.4035 ;
 END
 END vss.gds2158
 PIN vss.gds2159
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.39 26.2035 21.45 26.4035 ;
 END
 END vss.gds2159
 PIN vss.gds2160
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.726 26.2035 21.786 26.4035 ;
 END
 END vss.gds2160
 PIN vss.gds2161
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.894 26.2035 21.954 26.4035 ;
 END
 END vss.gds2161
 PIN vss.gds2162
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.062 26.2035 22.122 26.4035 ;
 END
 END vss.gds2162
 PIN vss.gds2163
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.398 26.2035 22.458 26.4035 ;
 END
 END vss.gds2163
 PIN vss.gds2164
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.566 26.2035 22.626 26.4035 ;
 END
 END vss.gds2164
 PIN vss.gds2165
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.734 26.2035 22.794 26.4035 ;
 END
 END vss.gds2165
 PIN vss.gds2166
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.07 26.2035 23.13 26.4035 ;
 END
 END vss.gds2166
 PIN vss.gds2167
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.238 26.2035 23.298 26.4035 ;
 END
 END vss.gds2167
 PIN vss.gds2168
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.406 26.2035 23.466 26.4035 ;
 END
 END vss.gds2168
 PIN vss.gds2169
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 27.092 24.726 27.292 ;
 END
 END vss.gds2169
 PIN vss.gds2170
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 27.092 22.962 27.292 ;
 END
 END vss.gds2170
 PIN vss.gds2171
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 27.092 22.29 27.292 ;
 END
 END vss.gds2171
 PIN vss.gds2172
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 27.092 21.618 27.292 ;
 END
 END vss.gds2172
 PIN vss.gds2173
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 27.092 20.946 27.292 ;
 END
 END vss.gds2173
 PIN vss.gds2174
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 27.092 23.634 27.292 ;
 END
 END vss.gds2174
 PIN vss.gds2175
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 23.912 25.52 23.968 25.72 ;
 RECT 23.912 26.78 23.968 26.98 ;
 RECT 23.912 28.04 23.968 28.24 ;
 RECT 23.744 27.1235 23.8 27.3235 ;
 END
 END vss.gds2175
 PIN vss.gds2176
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.202 26.2035 29.262 26.4035 ;
 END
 END vss.gds2176
 PIN vss.gds2177
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.034 26.2035 29.094 26.4035 ;
 END
 END vss.gds2177
 PIN vss.gds2178
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.866 26.2035 28.926 26.4035 ;
 END
 END vss.gds2178
 PIN vss.gds2179
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.53 26.2035 28.59 26.4035 ;
 END
 END vss.gds2179
 PIN vss.gds2180
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.362 26.2035 28.422 26.4035 ;
 END
 END vss.gds2180
 PIN vss.gds2181
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.194 26.2035 28.254 26.4035 ;
 END
 END vss.gds2181
 PIN vss.gds2182
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.858 26.2035 27.918 26.4035 ;
 END
 END vss.gds2182
 PIN vss.gds2183
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.69 26.2035 27.75 26.4035 ;
 END
 END vss.gds2183
 PIN vss.gds2184
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.522 26.2035 27.582 26.4035 ;
 END
 END vss.gds2184
 PIN vss.gds2185
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.186 26.2035 27.246 26.4035 ;
 END
 END vss.gds2185
 PIN vss.gds2186
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.018 26.2035 27.078 26.4035 ;
 END
 END vss.gds2186
 PIN vss.gds2187
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.85 26.2035 26.91 26.4035 ;
 END
 END vss.gds2187
 PIN vss.gds2188
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.514 26.2035 26.574 26.4035 ;
 END
 END vss.gds2188
 PIN vss.gds2189
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.346 26.2035 26.406 26.4035 ;
 END
 END vss.gds2189
 PIN vss.gds2190
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.178 26.2035 26.238 26.4035 ;
 END
 END vss.gds2190
 PIN vss.gds2191
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.842 26.2035 25.902 26.4035 ;
 END
 END vss.gds2191
 PIN vss.gds2192
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.674 26.2035 25.734 26.4035 ;
 END
 END vss.gds2192
 PIN vss.gds2193
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.506 26.2035 25.566 26.4035 ;
 END
 END vss.gds2193
 PIN vss.gds2194
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 26.9805 29.43 27.1805 ;
 END
 END vss.gds2194
 PIN vss.gds2195
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 27.092 28.758 27.292 ;
 END
 END vss.gds2195
 PIN vss.gds2196
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 27.092 28.086 27.292 ;
 END
 END vss.gds2196
 PIN vss.gds2197
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 27.092 27.414 27.292 ;
 END
 END vss.gds2197
 PIN vss.gds2198
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 27.092 26.742 27.292 ;
 END
 END vss.gds2198
 PIN vss.gds2199
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 27.092 26.07 27.292 ;
 END
 END vss.gds2199
 PIN vss.gds2200
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 27.092 25.398 27.292 ;
 END
 END vss.gds2200
 PIN vss.gds2201
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 26.568 30.11 26.768 ;
 END
 END vss.gds2201
 PIN vss.gds2202
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 27.1335 29.87 27.3335 ;
 END
 END vss.gds2202
 PIN vss.gds2203
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 27.247 29.642 27.447 ;
 END
 END vss.gds2203
 PIN vss.gds2204
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.876 28.67 29.932 28.87 ;
 RECT 29.876 26.068 29.932 26.268 ;
 RECT 30.212 28.67 30.268 28.87 ;
 RECT 30.212 26.068 30.268 26.268 ;
 RECT 29.54 28.67 29.596 28.87 ;
 RECT 29.54 26.098 29.596 26.298 ;
 RECT 29.708 28.67 29.764 28.87 ;
 RECT 29.708 26.098 29.764 26.298 ;
 RECT 30.044 28.67 30.1 28.87 ;
 RECT 30.044 26.068 30.1 26.268 ;
 END
 END vss.gds2204
 PIN vss.gds2205
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 28.382 30.95 28.582 ;
 END
 END vss.gds2205
 PIN vss.gds2206
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 28.422 31.922 28.622 ;
 END
 END vss.gds2206
 PIN vss.gds2207
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 25.902 31.922 26.102 ;
 END
 END vss.gds2207
 PIN vss.gds2208
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 27.162 31.922 27.362 ;
 END
 END vss.gds2208
 PIN vss.gds2209
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 25.862 30.95 26.062 ;
 END
 END vss.gds2209
 PIN vss.gds2210
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 27.99 32.47 28.19 ;
 END
 END vss.gds2210
 PIN vss.gds2211
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.038 25.987 35.078 26.187 ;
 END
 END vss.gds2211
 PIN vss.gds2212
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.314 27.777 30.37 27.977 ;
 END
 END vss.gds2212
 PIN vss.gds2213
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 27.877 33.198 28.077 ;
 END
 END vss.gds2213
 PIN vss.gds2214
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 26.617 33.198 26.817 ;
 END
 END vss.gds2214
 PIN vss.gds2215
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 27.247 32.894 27.447 ;
 END
 END vss.gds2215
 PIN vss.gds2216
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 27.247 32.214 27.447 ;
 END
 END vss.gds2216
 PIN vss.gds2217
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.49 27.5195 34.546 27.7195 ;
 END
 END vss.gds2217
 PIN vss.gds2218
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 27.092 30.71 27.292 ;
 END
 END vss.gds2218
 PIN vss.gds2219
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 26.4895 33.866 26.6895 ;
 END
 END vss.gds2219
 PIN vss.gds2220
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 27.122 30.95 27.322 ;
 END
 END vss.gds2220
 PIN vss.gds2221
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 27.2705 33.542 27.4705 ;
 END
 END vss.gds2221
 PIN vss.gds2222
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 27.9975 34.366 28.1975 ;
 END
 END vss.gds2222
 PIN vss.gds2223
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 27.247 31.55 27.447 ;
 END
 END vss.gds2223
 PIN vss.gds2224
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 27.1335 34.886 27.3335 ;
 END
 END vss.gds2224
 PIN vss.gds2225
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 27.0605 34.046 27.2605 ;
 END
 END vss.gds2225
 PIN vss.gds2226
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 32.648 27.544 32.704 27.744 ;
 RECT 32.9 27.547 32.956 27.747 ;
 RECT 33.572 28.58 33.628 28.733 ;
 RECT 31.052 28.56 31.108 28.733 ;
 RECT 31.22 28.533 31.276 28.733 ;
 RECT 32.816 28.577 32.872 28.742 ;
 RECT 32.648 28.577 32.704 28.742 ;
 RECT 31.892 28.577 31.948 28.742 ;
 RECT 31.724 28.577 31.78 28.742 ;
 RECT 31.388 27.893 31.444 28.093 ;
 RECT 31.22 27.893 31.276 28.093 ;
 RECT 30.716 28.027 30.772 28.227 ;
 RECT 32.648 26.284 32.704 26.484 ;
 RECT 32.9 26.287 32.956 26.487 ;
 RECT 33.572 27.32 33.628 27.473 ;
 RECT 31.052 27.3 31.108 27.473 ;
 RECT 31.22 27.273 31.276 27.473 ;
 RECT 32.816 27.317 32.872 27.482 ;
 RECT 32.648 27.317 32.704 27.482 ;
 RECT 31.892 27.317 31.948 27.482 ;
 RECT 31.724 27.317 31.78 27.482 ;
 RECT 33.572 26.06 33.628 26.213 ;
 RECT 31.052 26.04 31.108 26.213 ;
 RECT 31.22 26.013 31.276 26.213 ;
 RECT 32.816 26.057 32.872 26.222 ;
 RECT 32.648 26.057 32.704 26.222 ;
 RECT 31.892 26.057 31.948 26.222 ;
 RECT 31.724 26.057 31.78 26.222 ;
 RECT 32.06 28.103 32.116 28.303 ;
 RECT 32.48 28.103 32.536 28.303 ;
 RECT 31.388 26.633 31.444 26.833 ;
 RECT 31.22 26.633 31.276 26.833 ;
 RECT 32.06 26.843 32.116 27.043 ;
 RECT 32.48 26.843 32.536 27.043 ;
 RECT 33.404 25.6835 33.46 25.8835 ;
 RECT 32.06 25.583 32.116 25.783 ;
 RECT 32.48 25.583 32.536 25.783 ;
 RECT 30.716 25.507 30.772 25.707 ;
 RECT 30.716 26.767 30.772 26.967 ;
 RECT 33.404 26.9435 33.46 27.1435 ;
 RECT 33.908 26.6915 33.964 26.8915 ;
 RECT 30.548 26.079 30.604 26.279 ;
 RECT 33.908 27.9515 33.964 28.1515 ;
 RECT 33.404 28.2035 33.46 28.4035 ;
 RECT 32.228 26.2835 32.284 26.4835 ;
 RECT 30.38 28.67 30.436 28.87 ;
 RECT 30.38 26.017 30.436 26.217 ;
 RECT 34.916 28.67 34.972 28.87 ;
 RECT 34.916 26.098 34.972 26.298 ;
 RECT 34.748 28.67 34.804 28.87 ;
 RECT 34.748 26.1055 34.804 26.3055 ;
 RECT 34.58 28.67 34.636 28.87 ;
 RECT 34.58 26.098 34.636 26.298 ;
 RECT 34.412 28.67 34.468 28.87 ;
 RECT 34.412 26.098 34.468 26.298 ;
 RECT 34.244 28.67 34.3 28.87 ;
 RECT 34.244 26.098 34.3 26.298 ;
 RECT 35.084 28.67 35.14 28.87 ;
 RECT 35.084 26.098 35.14 26.298 ;
 RECT 34.076 26.213 34.132 26.413 ;
 END
 END vss.gds2226
 PIN vss.gds2227
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.122 26.2035 40.182 26.4035 ;
 END
 END vss.gds2227
 PIN vss.gds2228
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.754 26.2035 35.814 26.4035 ;
 END
 END vss.gds2228
 PIN vss.gds2229
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.09 26.2035 36.15 26.4035 ;
 END
 END vss.gds2229
 PIN vss.gds2230
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.258 26.2035 36.318 26.4035 ;
 END
 END vss.gds2230
 PIN vss.gds2231
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.426 26.2035 36.486 26.4035 ;
 END
 END vss.gds2231
 PIN vss.gds2232
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.762 26.2035 36.822 26.4035 ;
 END
 END vss.gds2232
 PIN vss.gds2233
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.93 26.2035 36.99 26.4035 ;
 END
 END vss.gds2233
 PIN vss.gds2234
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.098 26.2035 37.158 26.4035 ;
 END
 END vss.gds2234
 PIN vss.gds2235
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.434 26.2035 37.494 26.4035 ;
 END
 END vss.gds2235
 PIN vss.gds2236
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.602 26.2035 37.662 26.4035 ;
 END
 END vss.gds2236
 PIN vss.gds2237
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.77 26.2035 37.83 26.4035 ;
 END
 END vss.gds2237
 PIN vss.gds2238
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.106 26.2035 38.166 26.4035 ;
 END
 END vss.gds2238
 PIN vss.gds2239
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.274 26.2035 38.334 26.4035 ;
 END
 END vss.gds2239
 PIN vss.gds2240
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.442 26.2035 38.502 26.4035 ;
 END
 END vss.gds2240
 PIN vss.gds2241
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 27.092 37.998 27.292 ;
 END
 END vss.gds2241
 PIN vss.gds2242
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 27.092 37.326 27.292 ;
 END
 END vss.gds2242
 PIN vss.gds2243
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 27.092 38.67 27.292 ;
 END
 END vss.gds2243
 PIN vss.gds2244
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.778 26.2035 38.838 26.4035 ;
 END
 END vss.gds2244
 PIN vss.gds2245
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.946 26.2035 39.006 26.4035 ;
 END
 END vss.gds2245
 PIN vss.gds2246
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.114 26.2035 39.174 26.4035 ;
 END
 END vss.gds2246
 PIN vss.gds2247
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.45 26.2035 39.51 26.4035 ;
 END
 END vss.gds2247
 PIN vss.gds2248
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.618 26.2035 39.678 26.4035 ;
 END
 END vss.gds2248
 PIN vss.gds2249
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.786 26.2035 39.846 26.4035 ;
 END
 END vss.gds2249
 PIN vss.gds2250
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.586 26.2035 35.646 26.4035 ;
 END
 END vss.gds2250
 PIN vss.gds2251
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.418 26.2035 35.478 26.4035 ;
 END
 END vss.gds2251
 PIN vss.gds2252
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 27.092 36.654 27.292 ;
 END
 END vss.gds2252
 PIN vss.gds2253
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 27.092 39.342 27.292 ;
 END
 END vss.gds2253
 PIN vss.gds2254
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 27.092 40.014 27.292 ;
 END
 END vss.gds2254
 PIN vss.gds2255
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 26.9805 35.31 27.1805 ;
 END
 END vss.gds2255
 PIN vss.gds2256
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 27.092 35.982 27.292 ;
 END
 END vss.gds2256
 PIN vss.gds2257
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.91 26.2035 44.97 26.4035 ;
 END
 END vss.gds2257
 PIN vss.gds2258
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.742 26.2035 44.802 26.4035 ;
 END
 END vss.gds2258
 PIN vss.gds2259
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.574 26.2035 44.634 26.4035 ;
 END
 END vss.gds2259
 PIN vss.gds2260
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.238 26.2035 44.298 26.4035 ;
 END
 END vss.gds2260
 PIN vss.gds2261
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.07 26.2035 44.13 26.4035 ;
 END
 END vss.gds2261
 PIN vss.gds2262
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.902 26.2035 43.962 26.4035 ;
 END
 END vss.gds2262
 PIN vss.gds2263
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.566 26.2035 43.626 26.4035 ;
 END
 END vss.gds2263
 PIN vss.gds2264
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.398 26.2035 43.458 26.4035 ;
 END
 END vss.gds2264
 PIN vss.gds2265
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.23 26.2035 43.29 26.4035 ;
 END
 END vss.gds2265
 PIN vss.gds2266
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.894 26.2035 42.954 26.4035 ;
 END
 END vss.gds2266
 PIN vss.gds2267
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.726 26.2035 42.786 26.4035 ;
 END
 END vss.gds2267
 PIN vss.gds2268
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.558 26.2035 42.618 26.4035 ;
 END
 END vss.gds2268
 PIN vss.gds2269
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.222 26.2035 42.282 26.4035 ;
 END
 END vss.gds2269
 PIN vss.gds2270
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.054 26.2035 42.114 26.4035 ;
 END
 END vss.gds2270
 PIN vss.gds2271
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.886 26.2035 41.946 26.4035 ;
 END
 END vss.gds2271
 PIN vss.gds2272
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.55 26.2035 41.61 26.4035 ;
 END
 END vss.gds2272
 PIN vss.gds2273
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.382 26.2035 41.442 26.4035 ;
 END
 END vss.gds2273
 PIN vss.gds2274
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.214 26.2035 41.274 26.4035 ;
 END
 END vss.gds2274
 PIN vss.gds2275
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.29 26.2035 40.35 26.4035 ;
 END
 END vss.gds2275
 PIN vss.gds2276
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.458 26.2035 40.518 26.4035 ;
 END
 END vss.gds2276
 PIN vss.gds2277
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 27.092 45.138 27.292 ;
 END
 END vss.gds2277
 PIN vss.gds2278
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 27.092 44.466 27.292 ;
 END
 END vss.gds2278
 PIN vss.gds2279
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 27.092 43.794 27.292 ;
 END
 END vss.gds2279
 PIN vss.gds2280
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 27.092 43.122 27.292 ;
 END
 END vss.gds2280
 PIN vss.gds2281
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 27.092 42.45 27.292 ;
 END
 END vss.gds2281
 PIN vss.gds2282
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 27.092 41.778 27.292 ;
 END
 END vss.gds2282
 PIN vss.gds2283
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 27.092 40.686 27.292 ;
 END
 END vss.gds2283
 PIN vss.gds2284
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 40.964 26.78 41.02 26.98 ;
 RECT 40.964 25.52 41.02 25.72 ;
 RECT 40.964 28.04 41.02 28.24 ;
 RECT 40.796 27.1235 40.852 27.3235 ;
 END
 END vss.gds2284
 PIN vss.gds2285
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 28.382 48.002 28.582 ;
 END
 END vss.gds2285
 PIN vss.gds2286
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 28.422 48.974 28.622 ;
 END
 END vss.gds2286
 PIN vss.gds2287
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 25.902 48.974 26.102 ;
 END
 END vss.gds2287
 PIN vss.gds2288
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 27.162 48.974 27.362 ;
 END
 END vss.gds2288
 PIN vss.gds2289
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 25.862 48.002 26.062 ;
 END
 END vss.gds2289
 PIN vss.gds2290
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 27.122 48.002 27.322 ;
 END
 END vss.gds2290
 PIN vss.gds2291
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 27.99 49.522 28.19 ;
 END
 END vss.gds2291
 PIN vss.gds2292
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.366 27.777 47.422 27.977 ;
 END
 END vss.gds2292
 PIN vss.gds2293
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.254 26.2035 46.314 26.4035 ;
 END
 END vss.gds2293
 PIN vss.gds2294
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.086 26.2035 46.146 26.4035 ;
 END
 END vss.gds2294
 PIN vss.gds2295
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.918 26.2035 45.978 26.4035 ;
 END
 END vss.gds2295
 PIN vss.gds2296
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.582 26.2035 45.642 26.4035 ;
 END
 END vss.gds2296
 PIN vss.gds2297
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.414 26.2035 45.474 26.4035 ;
 END
 END vss.gds2297
 PIN vss.gds2298
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.246 26.2035 45.306 26.4035 ;
 END
 END vss.gds2298
 PIN vss.gds2299
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 27.092 45.81 27.292 ;
 END
 END vss.gds2299
 PIN vss.gds2300
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 26.9805 46.482 27.1805 ;
 END
 END vss.gds2300
 PIN vss.gds2301
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 26.568 47.162 26.768 ;
 END
 END vss.gds2301
 PIN vss.gds2302
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 27.877 50.25 28.077 ;
 END
 END vss.gds2302
 PIN vss.gds2303
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 26.617 50.25 26.817 ;
 END
 END vss.gds2303
 PIN vss.gds2304
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 27.1335 46.922 27.3335 ;
 END
 END vss.gds2304
 PIN vss.gds2305
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 27.247 46.694 27.447 ;
 END
 END vss.gds2305
 PIN vss.gds2306
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 27.092 47.762 27.292 ;
 END
 END vss.gds2306
 PIN vss.gds2307
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 27.247 49.266 27.447 ;
 END
 END vss.gds2307
 PIN vss.gds2308
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 27.247 48.602 27.447 ;
 END
 END vss.gds2308
 PIN vss.gds2309
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 27.247 49.946 27.447 ;
 END
 END vss.gds2309
 PIN vss.gds2310
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 48.104 28.56 48.16 28.733 ;
 RECT 48.272 28.533 48.328 28.733 ;
 RECT 49.868 28.577 49.924 28.742 ;
 RECT 49.7 28.577 49.756 28.742 ;
 RECT 48.944 28.577 49 28.742 ;
 RECT 48.776 28.577 48.832 28.742 ;
 RECT 49.7 27.544 49.756 27.744 ;
 RECT 49.952 27.547 50.008 27.747 ;
 RECT 48.104 27.3 48.16 27.473 ;
 RECT 48.272 27.273 48.328 27.473 ;
 RECT 49.868 27.317 49.924 27.482 ;
 RECT 49.7 27.317 49.756 27.482 ;
 RECT 48.944 27.317 49 27.482 ;
 RECT 48.776 27.317 48.832 27.482 ;
 RECT 48.44 27.893 48.496 28.093 ;
 RECT 48.272 27.893 48.328 28.093 ;
 RECT 47.768 28.027 47.824 28.227 ;
 RECT 48.104 26.04 48.16 26.213 ;
 RECT 48.272 26.013 48.328 26.213 ;
 RECT 49.868 26.057 49.924 26.222 ;
 RECT 49.7 26.057 49.756 26.222 ;
 RECT 48.944 26.057 49 26.222 ;
 RECT 48.776 26.057 48.832 26.222 ;
 RECT 49.7 26.284 49.756 26.484 ;
 RECT 49.952 26.287 50.008 26.487 ;
 RECT 49.112 28.103 49.168 28.303 ;
 RECT 49.532 28.103 49.588 28.303 ;
 RECT 49.112 25.583 49.168 25.783 ;
 RECT 49.112 26.843 49.168 27.043 ;
 RECT 49.532 26.843 49.588 27.043 ;
 RECT 48.44 26.633 48.496 26.833 ;
 RECT 48.272 26.633 48.328 26.833 ;
 RECT 47.768 26.767 47.824 26.967 ;
 RECT 47.768 25.507 47.824 25.707 ;
 RECT 49.532 25.583 49.588 25.783 ;
 RECT 47.6 26.079 47.656 26.279 ;
 RECT 46.928 28.67 46.984 28.87 ;
 RECT 46.928 26.068 46.984 26.268 ;
 RECT 46.592 28.67 46.648 28.87 ;
 RECT 46.592 26.098 46.648 26.298 ;
 RECT 47.432 28.67 47.488 28.87 ;
 RECT 47.432 26.017 47.488 26.217 ;
 RECT 46.76 28.67 46.816 28.87 ;
 RECT 46.76 26.098 46.816 26.298 ;
 RECT 49.28 26.2835 49.336 26.4835 ;
 RECT 47.264 28.67 47.32 28.87 ;
 RECT 47.264 26.068 47.32 26.268 ;
 RECT 47.096 28.67 47.152 28.87 ;
 RECT 47.096 26.068 47.152 26.268 ;
 END
 END vss.gds2310
 PIN vss.gds2311
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.638 26.2035 52.698 26.4035 ;
 END
 END vss.gds2311
 PIN vss.gds2312
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.806 26.2035 52.866 26.4035 ;
 END
 END vss.gds2312
 PIN vss.gds2313
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.142 26.2035 53.202 26.4035 ;
 END
 END vss.gds2313
 PIN vss.gds2314
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.31 26.2035 53.37 26.4035 ;
 END
 END vss.gds2314
 PIN vss.gds2315
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.478 26.2035 53.538 26.4035 ;
 END
 END vss.gds2315
 PIN vss.gds2316
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.814 26.2035 53.874 26.4035 ;
 END
 END vss.gds2316
 PIN vss.gds2317
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.982 26.2035 54.042 26.4035 ;
 END
 END vss.gds2317
 PIN vss.gds2318
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.15 26.2035 54.21 26.4035 ;
 END
 END vss.gds2318
 PIN vss.gds2319
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 27.092 54.378 27.292 ;
 END
 END vss.gds2319
 PIN vss.gds2320
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.486 26.2035 54.546 26.4035 ;
 END
 END vss.gds2320
 PIN vss.gds2321
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.654 26.2035 54.714 26.4035 ;
 END
 END vss.gds2321
 PIN vss.gds2322
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.822 26.2035 54.882 26.4035 ;
 END
 END vss.gds2322
 PIN vss.gds2323
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 27.092 55.05 27.292 ;
 END
 END vss.gds2323
 PIN vss.gds2324
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.158 26.2035 55.218 26.4035 ;
 END
 END vss.gds2324
 PIN vss.gds2325
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 26.4895 50.918 26.6895 ;
 END
 END vss.gds2325
 PIN vss.gds2326
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.542 27.5195 51.598 27.7195 ;
 END
 END vss.gds2326
 PIN vss.gds2327
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 27.092 53.706 27.292 ;
 END
 END vss.gds2327
 PIN vss.gds2328
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.47 26.2035 52.53 26.4035 ;
 END
 END vss.gds2328
 PIN vss.gds2329
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 27.9975 51.418 28.1975 ;
 END
 END vss.gds2329
 PIN vss.gds2330
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 27.092 53.034 27.292 ;
 END
 END vss.gds2330
 PIN vss.gds2331
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.09 25.987 52.13 26.187 ;
 END
 END vss.gds2331
 PIN vss.gds2332
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 27.1335 51.938 27.3335 ;
 END
 END vss.gds2332
 PIN vss.gds2333
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 27.2705 50.594 27.4705 ;
 END
 END vss.gds2333
 PIN vss.gds2334
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 26.9805 52.362 27.1805 ;
 END
 END vss.gds2334
 PIN vss.gds2335
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 27.0605 51.098 27.2605 ;
 END
 END vss.gds2335
 PIN vss.gds2336
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 50.624 28.58 50.68 28.733 ;
 RECT 50.624 27.32 50.68 27.473 ;
 RECT 50.624 26.06 50.68 26.213 ;
 RECT 50.456 25.6835 50.512 25.8835 ;
 RECT 50.96 26.6915 51.016 26.8915 ;
 RECT 50.456 26.9435 50.512 27.1435 ;
 RECT 50.96 27.9515 51.016 28.1515 ;
 RECT 50.456 28.2035 50.512 28.4035 ;
 RECT 51.968 28.67 52.024 28.87 ;
 RECT 51.968 26.098 52.024 26.298 ;
 RECT 51.8 28.67 51.856 28.87 ;
 RECT 51.8 26.1055 51.856 26.3055 ;
 RECT 51.632 28.67 51.688 28.87 ;
 RECT 51.632 26.098 51.688 26.298 ;
 RECT 51.464 28.67 51.52 28.87 ;
 RECT 51.464 26.098 51.52 26.298 ;
 RECT 51.296 28.67 51.352 28.87 ;
 RECT 51.296 26.098 51.352 26.298 ;
 RECT 51.128 26.213 51.184 26.413 ;
 RECT 52.136 28.67 52.192 28.87 ;
 RECT 52.136 26.098 52.192 26.298 ;
 END
 END vss.gds2336
 PIN vss.gds2337
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 27.092 60.174 27.292 ;
 END
 END vss.gds2337
 PIN vss.gds2338
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.946 26.2035 60.006 26.4035 ;
 END
 END vss.gds2338
 PIN vss.gds2339
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.778 26.2035 59.838 26.4035 ;
 END
 END vss.gds2339
 PIN vss.gds2340
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.61 26.2035 59.67 26.4035 ;
 END
 END vss.gds2340
 PIN vss.gds2341
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 27.092 59.502 27.292 ;
 END
 END vss.gds2341
 PIN vss.gds2342
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.274 26.2035 59.334 26.4035 ;
 END
 END vss.gds2342
 PIN vss.gds2343
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.106 26.2035 59.166 26.4035 ;
 END
 END vss.gds2343
 PIN vss.gds2344
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.938 26.2035 58.998 26.4035 ;
 END
 END vss.gds2344
 PIN vss.gds2345
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 27.092 58.83 27.292 ;
 END
 END vss.gds2345
 PIN vss.gds2346
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.602 26.2035 58.662 26.4035 ;
 END
 END vss.gds2346
 PIN vss.gds2347
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.434 26.2035 58.494 26.4035 ;
 END
 END vss.gds2347
 PIN vss.gds2348
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.266 26.2035 58.326 26.4035 ;
 END
 END vss.gds2348
 PIN vss.gds2349
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.326 26.2035 55.386 26.4035 ;
 END
 END vss.gds2349
 PIN vss.gds2350
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.494 26.2035 55.554 26.4035 ;
 END
 END vss.gds2350
 PIN vss.gds2351
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 27.092 55.722 27.292 ;
 END
 END vss.gds2351
 PIN vss.gds2352
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.83 26.2035 55.89 26.4035 ;
 END
 END vss.gds2352
 PIN vss.gds2353
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.998 26.2035 56.058 26.4035 ;
 END
 END vss.gds2353
 PIN vss.gds2354
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.166 26.2035 56.226 26.4035 ;
 END
 END vss.gds2354
 PIN vss.gds2355
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.502 26.2035 56.562 26.4035 ;
 END
 END vss.gds2355
 PIN vss.gds2356
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.67 26.2035 56.73 26.4035 ;
 END
 END vss.gds2356
 PIN vss.gds2357
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.838 26.2035 56.898 26.4035 ;
 END
 END vss.gds2357
 PIN vss.gds2358
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.342 26.2035 57.402 26.4035 ;
 END
 END vss.gds2358
 PIN vss.gds2359
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.51 26.2035 57.57 26.4035 ;
 END
 END vss.gds2359
 PIN vss.gds2360
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.174 26.2035 57.234 26.4035 ;
 END
 END vss.gds2360
 PIN vss.gds2361
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 27.092 56.394 27.292 ;
 END
 END vss.gds2361
 PIN vss.gds2362
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 27.092 57.738 27.292 ;
 END
 END vss.gds2362
 PIN vss.gds2363
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 27.092 57.066 27.292 ;
 END
 END vss.gds2363
 PIN vss.gds2364
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 58.016 25.52 58.072 25.72 ;
 RECT 58.016 26.78 58.072 26.98 ;
 RECT 58.016 28.04 58.072 28.24 ;
 RECT 57.848 27.1235 57.904 27.3235 ;
 END
 END vss.gds2364
 PIN vss.gds2365
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 28.382 65.054 28.582 ;
 END
 END vss.gds2365
 PIN vss.gds2366
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 25.862 65.054 26.062 ;
 END
 END vss.gds2366
 PIN vss.gds2367
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 27.122 65.054 27.322 ;
 END
 END vss.gds2367
 PIN vss.gds2368
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 26.568 64.214 26.768 ;
 END
 END vss.gds2368
 PIN vss.gds2369
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.418 27.777 64.474 27.977 ;
 END
 END vss.gds2369
 PIN vss.gds2370
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 26.9805 63.534 27.1805 ;
 END
 END vss.gds2370
 PIN vss.gds2371
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.306 26.2035 63.366 26.4035 ;
 END
 END vss.gds2371
 PIN vss.gds2372
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.138 26.2035 63.198 26.4035 ;
 END
 END vss.gds2372
 PIN vss.gds2373
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.97 26.2035 63.03 26.4035 ;
 END
 END vss.gds2373
 PIN vss.gds2374
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 27.092 62.862 27.292 ;
 END
 END vss.gds2374
 PIN vss.gds2375
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.634 26.2035 62.694 26.4035 ;
 END
 END vss.gds2375
 PIN vss.gds2376
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.466 26.2035 62.526 26.4035 ;
 END
 END vss.gds2376
 PIN vss.gds2377
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.298 26.2035 62.358 26.4035 ;
 END
 END vss.gds2377
 PIN vss.gds2378
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 27.092 62.19 27.292 ;
 END
 END vss.gds2378
 PIN vss.gds2379
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.962 26.2035 62.022 26.4035 ;
 END
 END vss.gds2379
 PIN vss.gds2380
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.794 26.2035 61.854 26.4035 ;
 END
 END vss.gds2380
 PIN vss.gds2381
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.626 26.2035 61.686 26.4035 ;
 END
 END vss.gds2381
 PIN vss.gds2382
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 27.092 61.518 27.292 ;
 END
 END vss.gds2382
 PIN vss.gds2383
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.29 26.2035 61.35 26.4035 ;
 END
 END vss.gds2383
 PIN vss.gds2384
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.122 26.2035 61.182 26.4035 ;
 END
 END vss.gds2384
 PIN vss.gds2385
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.954 26.2035 61.014 26.4035 ;
 END
 END vss.gds2385
 PIN vss.gds2386
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 27.092 60.846 27.292 ;
 END
 END vss.gds2386
 PIN vss.gds2387
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.618 26.2035 60.678 26.4035 ;
 END
 END vss.gds2387
 PIN vss.gds2388
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.45 26.2035 60.51 26.4035 ;
 END
 END vss.gds2388
 PIN vss.gds2389
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.282 26.2035 60.342 26.4035 ;
 END
 END vss.gds2389
 PIN vss.gds2390
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 27.1335 63.974 27.3335 ;
 END
 END vss.gds2390
 PIN vss.gds2391
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 27.247 63.746 27.447 ;
 END
 END vss.gds2391
 PIN vss.gds2392
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 27.092 64.814 27.292 ;
 END
 END vss.gds2392
 PIN vss.gds2393
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 65.156 28.56 65.212 28.733 ;
 RECT 65.156 27.3 65.212 27.473 ;
 RECT 65.156 26.04 65.212 26.213 ;
 RECT 64.82 28.027 64.876 28.227 ;
 RECT 64.82 26.767 64.876 26.967 ;
 RECT 64.82 25.507 64.876 25.707 ;
 RECT 64.652 26.079 64.708 26.279 ;
 RECT 63.98 28.67 64.036 28.87 ;
 RECT 63.98 26.068 64.036 26.268 ;
 RECT 64.484 28.67 64.54 28.87 ;
 RECT 64.484 26.017 64.54 26.217 ;
 RECT 63.812 28.67 63.868 28.87 ;
 RECT 63.812 26.098 63.868 26.298 ;
 RECT 64.316 28.67 64.372 28.87 ;
 RECT 64.316 26.068 64.372 26.268 ;
 RECT 64.148 28.67 64.204 28.87 ;
 RECT 64.148 26.068 64.204 26.268 ;
 RECT 63.644 28.67 63.7 28.87 ;
 RECT 63.644 26.098 63.7 26.298 ;
 END
 END vss.gds2393
 PIN vss.gds2394
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 28.422 66.026 28.622 ;
 END
 END vss.gds2394
 PIN vss.gds2395
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 25.902 66.026 26.102 ;
 END
 END vss.gds2395
 PIN vss.gds2396
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 27.162 66.026 27.362 ;
 END
 END vss.gds2396
 PIN vss.gds2397
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 27.247 66.318 27.447 ;
 END
 END vss.gds2397
 PIN vss.gds2398
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 27.99 66.574 28.19 ;
 END
 END vss.gds2398
 PIN vss.gds2399
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.142 25.987 69.182 26.187 ;
 END
 END vss.gds2399
 PIN vss.gds2400
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 27.877 67.302 28.077 ;
 END
 END vss.gds2400
 PIN vss.gds2401
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.69 26.2035 69.75 26.4035 ;
 END
 END vss.gds2401
 PIN vss.gds2402
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.858 26.2035 69.918 26.4035 ;
 END
 END vss.gds2402
 PIN vss.gds2403
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 27.092 70.086 27.292 ;
 END
 END vss.gds2403
 PIN vss.gds2404
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.194 26.2035 70.254 26.4035 ;
 END
 END vss.gds2404
 PIN vss.gds2405
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.594 27.5195 68.65 27.7195 ;
 END
 END vss.gds2405
 PIN vss.gds2406
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 26.4895 67.97 26.6895 ;
 END
 END vss.gds2406
 PIN vss.gds2407
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 26.617 67.302 26.817 ;
 END
 END vss.gds2407
 PIN vss.gds2408
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.522 26.2035 69.582 26.4035 ;
 END
 END vss.gds2408
 PIN vss.gds2409
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 27.0605 68.15 27.2605 ;
 END
 END vss.gds2409
 PIN vss.gds2410
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 27.9975 68.47 28.1975 ;
 END
 END vss.gds2410
 PIN vss.gds2411
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 27.2705 67.646 27.4705 ;
 END
 END vss.gds2411
 PIN vss.gds2412
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 27.247 65.654 27.447 ;
 END
 END vss.gds2412
 PIN vss.gds2413
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 27.247 66.998 27.447 ;
 END
 END vss.gds2413
 PIN vss.gds2414
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 27.1335 68.99 27.3335 ;
 END
 END vss.gds2414
 PIN vss.gds2415
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 26.9805 69.414 27.1805 ;
 END
 END vss.gds2415
 PIN vss.gds2416
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 66.752 27.544 66.808 27.744 ;
 RECT 67.004 27.547 67.06 27.747 ;
 RECT 67.676 28.58 67.732 28.733 ;
 RECT 65.324 28.533 65.38 28.733 ;
 RECT 66.92 28.577 66.976 28.742 ;
 RECT 66.752 28.577 66.808 28.742 ;
 RECT 65.996 28.577 66.052 28.742 ;
 RECT 65.828 28.577 65.884 28.742 ;
 RECT 67.676 27.32 67.732 27.473 ;
 RECT 65.324 27.273 65.38 27.473 ;
 RECT 66.92 27.317 66.976 27.482 ;
 RECT 66.752 27.317 66.808 27.482 ;
 RECT 65.996 27.317 66.052 27.482 ;
 RECT 65.828 27.317 65.884 27.482 ;
 RECT 67.676 26.06 67.732 26.213 ;
 RECT 65.324 26.013 65.38 26.213 ;
 RECT 66.92 26.057 66.976 26.222 ;
 RECT 66.752 26.057 66.808 26.222 ;
 RECT 65.996 26.057 66.052 26.222 ;
 RECT 65.828 26.057 65.884 26.222 ;
 RECT 65.492 27.893 65.548 28.093 ;
 RECT 65.324 27.893 65.38 28.093 ;
 RECT 66.752 26.284 66.808 26.484 ;
 RECT 67.004 26.287 67.06 26.487 ;
 RECT 66.164 28.103 66.22 28.303 ;
 RECT 66.584 28.103 66.64 28.303 ;
 RECT 66.164 26.843 66.22 27.043 ;
 RECT 66.584 26.843 66.64 27.043 ;
 RECT 65.492 26.633 65.548 26.833 ;
 RECT 65.324 26.633 65.38 26.833 ;
 RECT 67.508 26.9435 67.564 27.1435 ;
 RECT 68.012 26.6915 68.068 26.8915 ;
 RECT 67.508 25.6835 67.564 25.8835 ;
 RECT 66.164 25.583 66.22 25.783 ;
 RECT 66.584 25.583 66.64 25.783 ;
 RECT 68.012 27.9515 68.068 28.1515 ;
 RECT 67.508 28.2035 67.564 28.4035 ;
 RECT 66.332 26.2835 66.388 26.4835 ;
 RECT 69.02 28.67 69.076 28.87 ;
 RECT 69.02 26.098 69.076 26.298 ;
 RECT 68.852 28.67 68.908 28.87 ;
 RECT 68.852 26.1055 68.908 26.3055 ;
 RECT 68.684 28.67 68.74 28.87 ;
 RECT 68.684 26.098 68.74 26.298 ;
 RECT 68.516 28.67 68.572 28.87 ;
 RECT 68.516 26.098 68.572 26.298 ;
 RECT 68.348 28.67 68.404 28.87 ;
 RECT 68.348 26.098 68.404 26.298 ;
 RECT 69.188 28.67 69.244 28.87 ;
 RECT 69.188 26.098 69.244 26.298 ;
 RECT 68.18 26.213 68.236 26.413 ;
 END
 END vss.gds2416
 PIN vss.gds2417
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.362 26.2035 70.422 26.4035 ;
 END
 END vss.gds2417
 PIN vss.gds2418
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.53 26.2035 70.59 26.4035 ;
 END
 END vss.gds2418
 PIN vss.gds2419
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.866 26.2035 70.926 26.4035 ;
 END
 END vss.gds2419
 PIN vss.gds2420
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.034 26.2035 71.094 26.4035 ;
 END
 END vss.gds2420
 PIN vss.gds2421
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.202 26.2035 71.262 26.4035 ;
 END
 END vss.gds2421
 PIN vss.gds2422
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 27.092 71.43 27.292 ;
 END
 END vss.gds2422
 PIN vss.gds2423
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.538 26.2035 71.598 26.4035 ;
 END
 END vss.gds2423
 PIN vss.gds2424
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.706 26.2035 71.766 26.4035 ;
 END
 END vss.gds2424
 PIN vss.gds2425
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.874 26.2035 71.934 26.4035 ;
 END
 END vss.gds2425
 PIN vss.gds2426
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 27.092 72.102 27.292 ;
 END
 END vss.gds2426
 PIN vss.gds2427
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.21 26.2035 72.27 26.4035 ;
 END
 END vss.gds2427
 PIN vss.gds2428
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.378 26.2035 72.438 26.4035 ;
 END
 END vss.gds2428
 PIN vss.gds2429
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.546 26.2035 72.606 26.4035 ;
 END
 END vss.gds2429
 PIN vss.gds2430
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 27.092 72.774 27.292 ;
 END
 END vss.gds2430
 PIN vss.gds2431
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.882 26.2035 72.942 26.4035 ;
 END
 END vss.gds2431
 PIN vss.gds2432
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.05 26.2035 73.11 26.4035 ;
 END
 END vss.gds2432
 PIN vss.gds2433
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.554 26.2035 73.614 26.4035 ;
 END
 END vss.gds2433
 PIN vss.gds2434
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.722 26.2035 73.782 26.4035 ;
 END
 END vss.gds2434
 PIN vss.gds2435
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.89 26.2035 73.95 26.4035 ;
 END
 END vss.gds2435
 PIN vss.gds2436
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.226 26.2035 74.286 26.4035 ;
 END
 END vss.gds2436
 PIN vss.gds2437
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.394 26.2035 74.454 26.4035 ;
 END
 END vss.gds2437
 PIN vss.gds2438
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.218 26.2035 73.278 26.4035 ;
 END
 END vss.gds2438
 PIN vss.gds2439
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.562 26.2035 74.622 26.4035 ;
 END
 END vss.gds2439
 PIN vss.gds2440
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 27.092 70.758 27.292 ;
 END
 END vss.gds2440
 PIN vss.gds2441
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 27.092 74.118 27.292 ;
 END
 END vss.gds2441
 PIN vss.gds2442
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 27.092 74.79 27.292 ;
 END
 END vss.gds2442
 PIN vss.gds2443
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 27.092 73.446 27.292 ;
 END
 END vss.gds2443
 PIN vccdgt_1p0
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 4.979 0.654 5.179 ;
 END
 END vccdgt_1p0
 PIN vccdgt_1p0.gds1
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 3.719 0.654 3.919 ;
 END
 END vccdgt_1p0.gds1
 PIN vccdgt_1p0.gds2
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 2.459 0.654 2.659 ;
 END
 END vccdgt_1p0.gds2
 PIN vccdgt_1p0.gds3
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 1.199 0.654 1.399 ;
 END
 END vccdgt_1p0.gds3
 PIN vccdgt_1p0.gds4
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.454 2.978 0.494 3.178 ;
 END
 END vccdgt_1p0.gds4
 PIN vccdgt_1p0.gds5
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.742 3.0505 0.788 3.2505 ;
 END
 END vccdgt_1p0.gds5
 PIN vccdgt_1p0.gds6
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.114 3.003 1.154 3.203 ;
 END
 END vccdgt_1p0.gds6
 PIN vccdgt_1p0.gds7
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.566 2.903 1.622 3.103 ;
 END
 END vccdgt_1p0.gds7
 PIN vccdgt_1p0.gds8
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.166 2.966 3.206 3.166 ;
 END
 END vccdgt_1p0.gds8
 PIN vccdgt_1p0.gds9
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.966 2.9665 1.026 3.1665 ;
 END
 END vccdgt_1p0.gds9
 PIN vccdgt_1p0.gds10
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.986 3.0425 2.042 3.2425 ;
 END
 END vccdgt_1p0.gds10
 PIN vccdgt_1p0.gds11
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.326 3.0145 2.382 3.2145 ;
 END
 END vccdgt_1p0.gds11
 PIN vccdgt_1p0.gds12
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.806 3.052 1.882 3.252 ;
 END
 END vccdgt_1p0.gds12
 PIN vccdgt_1p0.gds13
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.646 2.9745 2.722 3.1745 ;
 END
 END vccdgt_1p0.gds13
 PIN vccdgt_1p0.gds14
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.634 3.139 4.674 3.339 ;
 END
 END vccdgt_1p0.gds14
 PIN vccdgt_1p0.gds15
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.098 2.9955 5.138 3.1955 ;
 END
 END vccdgt_1p0.gds15
 PIN vccdgt_1p0.gds16
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.478 2.98 3.538 3.18 ;
 END
 END vccdgt_1p0.gds16
 PIN vccdgt_1p0.gds17
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.69 3.059 3.73 3.259 ;
 END
 END vccdgt_1p0.gds17
 PIN vccdgt_1p0.gds18
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.882 3.0725 3.922 3.2725 ;
 END
 END vccdgt_1p0.gds18
 PIN vccdgt_1p0.gds19
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.362 3.058 4.418 3.258 ;
 END
 END vccdgt_1p0.gds19
 PIN vccdgt_1p0.gds20
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.09 3.0505 4.13 3.2505 ;
 END
 END vccdgt_1p0.gds20
 PIN vccdgt_1p0.gds21
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.906 3.082 4.946 3.282 ;
 END
 END vccdgt_1p0.gds21
 PIN vccdgt_1p0.gds22
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.762 2.978 4.818 3.178 ;
 END
 END vccdgt_1p0.gds22
 PIN vccdgt_1p0.gds23
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.486 3.058 2.542 3.258 ;
 END
 END vccdgt_1p0.gds23
 PIN vccdgt_1p0.gds24
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 1.232 1.476 1.288 1.676 ;
 RECT 1.568 1.491 1.624 1.691 ;
 RECT 1.82 1.491 1.876 1.691 ;
 RECT 2.072 1.605 2.128 1.785 ;
 RECT 2.996 1.603 3.052 1.785 ;
 RECT 3.164 1.603 3.22 1.779 ;
 RECT 2.492 1.1045 2.548 1.3045 ;
 RECT 1.232 2.736 1.288 2.936 ;
 RECT 1.568 2.751 1.624 2.951 ;
 RECT 1.82 2.751 1.876 2.951 ;
 RECT 2.072 2.865 2.128 3.045 ;
 RECT 2.996 2.863 3.052 3.045 ;
 RECT 3.164 2.863 3.22 3.039 ;
 RECT 2.492 2.3645 2.548 2.5645 ;
 RECT 1.232 3.996 1.288 4.196 ;
 RECT 1.568 4.011 1.624 4.211 ;
 RECT 1.82 4.011 1.876 4.211 ;
 RECT 2.072 4.125 2.128 4.305 ;
 RECT 2.996 4.123 3.052 4.305 ;
 RECT 3.164 4.123 3.22 4.299 ;
 RECT 2.492 3.6245 2.548 3.8245 ;
 RECT 1.232 5.256 1.288 5.456 ;
 RECT 1.568 5.271 1.624 5.471 ;
 RECT 1.82 5.271 1.876 5.471 ;
 RECT 2.072 5.385 2.128 5.565 ;
 RECT 2.996 5.383 3.052 5.565 ;
 RECT 3.164 5.383 3.22 5.559 ;
 RECT 2.492 4.8845 2.548 5.0845 ;
 RECT 0.812 1.509 0.868 1.709 ;
 RECT 0.644 1.509 0.7 1.709 ;
 RECT 0.98 1.509 1.036 1.709 ;
 RECT 0.812 2.769 0.868 2.969 ;
 RECT 0.644 2.769 0.7 2.969 ;
 RECT 0.98 2.769 1.036 2.969 ;
 RECT 0.812 4.029 0.868 4.229 ;
 RECT 0.644 4.029 0.7 4.229 ;
 RECT 0.98 4.029 1.036 4.229 ;
 RECT 0.812 5.289 0.868 5.489 ;
 RECT 0.644 5.289 0.7 5.489 ;
 RECT 0.98 5.289 1.036 5.489 ;
 RECT 4.088 4.8335 4.144 5.0335 ;
 RECT 4.676 4.8335 4.732 5.0335 ;
 RECT 4.424 4.8335 4.48 5.0335 ;
 RECT 5.012 4.8335 5.068 5.0335 ;
 RECT 4.844 4.8335 4.9 5.0335 ;
 RECT 4.088 3.5735 4.144 3.7735 ;
 RECT 4.676 3.5735 4.732 3.7735 ;
 RECT 4.424 3.5735 4.48 3.7735 ;
 RECT 5.012 3.5735 5.068 3.7735 ;
 RECT 4.844 3.5735 4.9 3.7735 ;
 RECT 4.088 2.3135 4.144 2.5135 ;
 RECT 4.676 2.3135 4.732 2.5135 ;
 RECT 4.424 2.3135 4.48 2.5135 ;
 RECT 5.012 2.3135 5.068 2.5135 ;
 RECT 4.844 2.3135 4.9 2.5135 ;
 RECT 4.088 1.0535 4.144 1.2535 ;
 RECT 4.676 1.0535 4.732 1.2535 ;
 RECT 4.424 1.0535 4.48 1.2535 ;
 RECT 5.012 1.0535 5.068 1.2535 ;
 RECT 4.844 1.0535 4.9 1.2535 ;
 END
 END vccdgt_1p0.gds24
 PIN vccdgt_1p0.gds25
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.33 3.209 6.37 3.409 ;
 END
 END vccdgt_1p0.gds25
 PIN vccdgt_1p0.gds26
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.498 2.98 5.538 3.18 ;
 END
 END vccdgt_1p0.gds26
 PIN vccdgt_1p0.gds27
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.862 3.0725 6.918 3.2725 ;
 END
 END vccdgt_1p0.gds27
 PIN vccdgt_1p0.gds28
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.074 3.082 6.114 3.282 ;
 END
 END vccdgt_1p0.gds28
 PIN vccdgt_1p0.gds29
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.306 3.0725 5.346 3.2725 ;
 END
 END vccdgt_1p0.gds29
 PIN vccdgt_1p0.gds30
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.818 3.0505 5.858 3.2505 ;
 END
 END vccdgt_1p0.gds30
 PIN vccdgt_1p0.gds31
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.626 2.951 5.666 3.151 ;
 END
 END vccdgt_1p0.gds31
 PIN vccdgt_1p0.gds32
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.202 3.0595 6.242 3.2595 ;
 END
 END vccdgt_1p0.gds32
 PIN vccdgt_1p0.gds33
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.67 2.999 6.71 3.199 ;
 END
 END vccdgt_1p0.gds33
 PIN vccdgt_1p0.gds34
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.348 4.8845 5.404 5.0845 ;
 RECT 6.02 4.8335 6.076 5.0335 ;
 RECT 5.684 4.9125 5.74 5.1125 ;
 RECT 6.356 4.9125 6.412 5.1125 ;
 RECT 5.348 3.6245 5.404 3.8245 ;
 RECT 6.02 3.5735 6.076 3.7735 ;
 RECT 5.684 3.6525 5.74 3.8525 ;
 RECT 6.356 3.6525 6.412 3.8525 ;
 RECT 5.348 2.3645 5.404 2.5645 ;
 RECT 6.02 2.3135 6.076 2.5135 ;
 RECT 5.684 2.3925 5.74 2.5925 ;
 RECT 6.356 2.3925 6.412 2.5925 ;
 RECT 5.348 1.1045 5.404 1.3045 ;
 RECT 6.02 1.0535 6.076 1.2535 ;
 RECT 5.684 1.1325 5.74 1.3325 ;
 RECT 6.356 1.1325 6.412 1.3325 ;
 END
 END vccdgt_1p0.gds34
 PIN vccdgt_1p0.gds35
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.522 3.1075 14.578 3.3075 ;
 END
 END vccdgt_1p0.gds35
 PIN vccdgt_1p0.gds36
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.342 2.8695 13.398 3.0695 ;
 END
 END vccdgt_1p0.gds36
 PIN vccdgt_1p0.gds37
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.186 3.1075 15.226 3.3075 ;
 END
 END vccdgt_1p0.gds37
 PIN vccdgt_1p0.gds38
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.502 2.82 13.558 3.02 ;
 END
 END vccdgt_1p0.gds38
 PIN vccdgt_1p0.gds39
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.182 3.25 14.238 3.45 ;
 END
 END vccdgt_1p0.gds39
 PIN vccdgt_1p0.gds40
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.766 3.054 14.806 3.254 ;
 END
 END vccdgt_1p0.gds40
 PIN vccdgt_1p0.gds41
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.678 3.0175 12.718 3.2175 ;
 END
 END vccdgt_1p0.gds41
 PIN vccdgt_1p0.gds42
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.162 2.9115 13.238 3.1115 ;
 END
 END vccdgt_1p0.gds42
 PIN vccdgt_1p0.gds43
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.002 3.25 14.078 3.45 ;
 END
 END vccdgt_1p0.gds43
 PIN vccdgt_1p0.gds44
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.958 3.3775 14.998 3.5775 ;
 END
 END vccdgt_1p0.gds44
 PIN vccdgt_1p0.gds45
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.402 2.9745 12.462 3.1745 ;
 END
 END vccdgt_1p0.gds45
 PIN vccdgt_1p0.gds46
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 14.756 1.013 14.812 1.213 ;
 RECT 14.756 2.273 14.812 2.473 ;
 RECT 14.756 3.533 14.812 3.733 ;
 RECT 14.756 4.793 14.812 4.993 ;
 RECT 14 4.676 14.056 4.876 ;
 RECT 14 0.896 14.056 1.096 ;
 RECT 14 2.156 14.056 2.356 ;
 RECT 14 3.416 14.056 3.616 ;
 RECT 14.924 4.36 14.98 4.56 ;
 RECT 14.588 4.793 14.644 4.993 ;
 RECT 14.42 4.78 14.476 4.98 ;
 RECT 14.924 3.1 14.98 3.3 ;
 RECT 14.588 3.533 14.644 3.733 ;
 RECT 14.42 3.52 14.476 3.72 ;
 RECT 14.924 1.84 14.98 2.04 ;
 RECT 14.588 2.273 14.644 2.473 ;
 RECT 14.42 2.26 14.476 2.46 ;
 RECT 14.924 0.58 14.98 0.78 ;
 RECT 14.588 1.013 14.644 1.213 ;
 RECT 14.42 1 14.476 1.2 ;
 END
 END vccdgt_1p0.gds46
 PIN vccdgt_1p0.gds47
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 4.042 16.57 4.242 ;
 END
 END vccdgt_1p0.gds47
 PIN vccdgt_1p0.gds48
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 2.782 16.57 2.982 ;
 END
 END vccdgt_1p0.gds48
 PIN vccdgt_1p0.gds49
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.018 2.862 17.074 3.062 ;
 END
 END vccdgt_1p0.gds49
 PIN vccdgt_1p0.gds50
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.838 2.8695 16.894 3.0695 ;
 END
 END vccdgt_1p0.gds50
 PIN vccdgt_1p0.gds51
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 5.302 16.57 5.502 ;
 END
 END vccdgt_1p0.gds51
 PIN vccdgt_1p0.gds52
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.866 3.1075 15.926 3.3075 ;
 END
 END vccdgt_1p0.gds52
 PIN vccdgt_1p0.gds53
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 1.522 16.57 1.722 ;
 END
 END vccdgt_1p0.gds53
 PIN vccdgt_1p0.gds54
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.03 3.265 16.076 3.465 ;
 END
 END vccdgt_1p0.gds54
 PIN vccdgt_1p0.gds55
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.314 3.054 15.354 3.254 ;
 END
 END vccdgt_1p0.gds55
 PIN vccdgt_1p0.gds56
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.338 2.8695 17.414 3.0695 ;
 END
 END vccdgt_1p0.gds56
 PIN vccdgt_1p0.gds57
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.522 3.0365 15.582 3.2365 ;
 END
 END vccdgt_1p0.gds57
 PIN vccdgt_1p0.gds58
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.598 3.0505 17.654 3.2505 ;
 END
 END vccdgt_1p0.gds58
 PIN vccdgt_1p0.gds59
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.674 2.8695 16.734 3.0695 ;
 END
 END vccdgt_1p0.gds59
 PIN vccdgt_1p0.gds60
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.858 3.016 17.898 3.216 ;
 END
 END vccdgt_1p0.gds60
 PIN vccdgt_1p0.gds61
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.114 2.9745 18.174 3.1745 ;
 END
 END vccdgt_1p0.gds61
 PIN vccdgt_1p0.gds62
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.178 3.016 17.234 3.216 ;
 END
 END vccdgt_1p0.gds62
 PIN vccdgt_1p0.gds63
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 15.932 1.076 15.988 1.276 ;
 RECT 16.1 2.273 16.156 2.473 ;
 RECT 15.932 4.856 15.988 5.056 ;
 RECT 15.764 4.436 15.82 4.636 ;
 RECT 15.512 4.688 15.568 4.888 ;
 RECT 15.26 4.775 15.316 4.975 ;
 RECT 16.1 4.793 16.156 4.993 ;
 RECT 15.764 3.176 15.82 3.376 ;
 RECT 15.512 3.428 15.568 3.628 ;
 RECT 15.932 3.596 15.988 3.796 ;
 RECT 16.1 3.533 16.156 3.733 ;
 RECT 15.26 3.515 15.316 3.715 ;
 RECT 15.764 1.916 15.82 2.116 ;
 RECT 15.512 2.168 15.568 2.368 ;
 RECT 15.932 2.336 15.988 2.536 ;
 RECT 15.26 2.255 15.316 2.455 ;
 RECT 15.764 0.656 15.82 0.856 ;
 RECT 15.512 0.908 15.568 1.108 ;
 RECT 15.26 0.995 15.316 1.195 ;
 RECT 16.1 1.013 16.156 1.213 ;
 END
 END vccdgt_1p0.gds63
 PIN vccdgt_1p0.gds64
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.93 2.978 23.97 3.178 ;
 END
 END vccdgt_1p0.gds64
 PIN vccdgt_1p0.gds65
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.658 2.979 23.698 3.179 ;
 END
 END vccdgt_1p0.gds65
 PIN vccdgt_1p0.gds66
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.214 2.9115 30.29 3.1115 ;
 END
 END vccdgt_1p0.gds66
 PIN vccdgt_1p0.gds67
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.73 3.0175 29.77 3.2175 ;
 END
 END vccdgt_1p0.gds67
 PIN vccdgt_1p0.gds68
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.454 2.9745 29.514 3.1745 ;
 END
 END vccdgt_1p0.gds68
 PIN vccdgt_1p0.gds69
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 5.302 33.622 5.502 ;
 END
 END vccdgt_1p0.gds69
 PIN vccdgt_1p0.gds70
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 4.042 33.622 4.242 ;
 END
 END vccdgt_1p0.gds70
 PIN vccdgt_1p0.gds71
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 2.782 33.622 2.982 ;
 END
 END vccdgt_1p0.gds71
 PIN vccdgt_1p0.gds72
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 1.522 33.622 1.722 ;
 END
 END vccdgt_1p0.gds72
 PIN vccdgt_1p0.gds73
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.07 2.862 34.126 3.062 ;
 END
 END vccdgt_1p0.gds73
 PIN vccdgt_1p0.gds74
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.89 2.8695 33.946 3.0695 ;
 END
 END vccdgt_1p0.gds74
 PIN vccdgt_1p0.gds75
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.918 3.1075 32.978 3.3075 ;
 END
 END vccdgt_1p0.gds75
 PIN vccdgt_1p0.gds76
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.574 3.1075 31.63 3.3075 ;
 END
 END vccdgt_1p0.gds76
 PIN vccdgt_1p0.gds77
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.394 2.8695 30.45 3.0695 ;
 END
 END vccdgt_1p0.gds77
 PIN vccdgt_1p0.gds78
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.39 2.8695 34.466 3.0695 ;
 END
 END vccdgt_1p0.gds78
 PIN vccdgt_1p0.gds79
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.238 3.054 32.278 3.254 ;
 END
 END vccdgt_1p0.gds79
 PIN vccdgt_1p0.gds80
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.818 3.054 31.858 3.254 ;
 END
 END vccdgt_1p0.gds80
 PIN vccdgt_1p0.gds81
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.234 3.25 31.29 3.45 ;
 END
 END vccdgt_1p0.gds81
 PIN vccdgt_1p0.gds82
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.082 3.265 33.128 3.465 ;
 END
 END vccdgt_1p0.gds82
 PIN vccdgt_1p0.gds83
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.366 3.1075 32.406 3.3075 ;
 END
 END vccdgt_1p0.gds83
 PIN vccdgt_1p0.gds84
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.01 3.3775 32.05 3.5775 ;
 END
 END vccdgt_1p0.gds84
 PIN vccdgt_1p0.gds85
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.166 2.9745 35.226 3.1745 ;
 END
 END vccdgt_1p0.gds85
 PIN vccdgt_1p0.gds86
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.91 3.016 34.95 3.216 ;
 END
 END vccdgt_1p0.gds86
 PIN vccdgt_1p0.gds87
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.054 3.25 31.13 3.45 ;
 END
 END vccdgt_1p0.gds87
 PIN vccdgt_1p0.gds88
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.554 2.82 30.61 3.02 ;
 END
 END vccdgt_1p0.gds88
 PIN vccdgt_1p0.gds89
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.23 3.016 34.286 3.216 ;
 END
 END vccdgt_1p0.gds89
 PIN vccdgt_1p0.gds90
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.65 3.0505 34.706 3.2505 ;
 END
 END vccdgt_1p0.gds90
 PIN vccdgt_1p0.gds91
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.574 3.0365 32.634 3.2365 ;
 END
 END vccdgt_1p0.gds91
 PIN vccdgt_1p0.gds92
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.726 2.8695 33.786 3.0695 ;
 END
 END vccdgt_1p0.gds92
 PIN vccdgt_1p0.gds93
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 31.808 1.013 31.864 1.213 ;
 RECT 32.984 1.076 33.04 1.276 ;
 RECT 33.152 2.273 33.208 2.473 ;
 RECT 31.808 2.273 31.864 2.473 ;
 RECT 31.808 3.533 31.864 3.733 ;
 RECT 33.152 4.793 33.208 4.993 ;
 RECT 31.808 4.793 31.864 4.993 ;
 RECT 31.052 0.896 31.108 1.096 ;
 RECT 31.052 2.156 31.108 2.356 ;
 RECT 31.052 3.416 31.108 3.616 ;
 RECT 31.052 4.676 31.108 4.876 ;
 RECT 31.976 4.36 32.032 4.56 ;
 RECT 32.816 4.436 32.872 4.636 ;
 RECT 32.564 4.688 32.62 4.888 ;
 RECT 32.984 4.856 33.04 5.056 ;
 RECT 32.312 4.775 32.368 4.975 ;
 RECT 31.64 4.793 31.696 4.993 ;
 RECT 31.472 4.78 31.528 4.98 ;
 RECT 31.976 3.1 32.032 3.3 ;
 RECT 32.816 3.176 32.872 3.376 ;
 RECT 32.564 3.428 32.62 3.628 ;
 RECT 32.984 3.596 33.04 3.796 ;
 RECT 33.152 3.533 33.208 3.733 ;
 RECT 31.64 3.533 31.696 3.733 ;
 RECT 31.472 3.52 31.528 3.72 ;
 RECT 32.312 3.515 32.368 3.715 ;
 RECT 31.976 1.84 32.032 2.04 ;
 RECT 32.816 1.916 32.872 2.116 ;
 RECT 32.564 2.168 32.62 2.368 ;
 RECT 32.984 2.336 33.04 2.536 ;
 RECT 32.312 2.255 32.368 2.455 ;
 RECT 31.64 2.273 31.696 2.473 ;
 RECT 31.472 2.26 31.528 2.46 ;
 RECT 31.976 0.58 32.032 0.78 ;
 RECT 32.816 0.656 32.872 0.856 ;
 RECT 32.564 0.908 32.62 1.108 ;
 RECT 32.312 0.995 32.368 1.195 ;
 RECT 31.64 1.013 31.696 1.213 ;
 RECT 33.152 1.013 33.208 1.213 ;
 RECT 31.472 1 31.528 1.2 ;
 END
 END vccdgt_1p0.gds93
 PIN vccdgt_1p0.gds94
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.982 2.978 41.022 3.178 ;
 END
 END vccdgt_1p0.gds94
 PIN vccdgt_1p0.gds95
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.71 2.979 40.75 3.179 ;
 END
 END vccdgt_1p0.gds95
 PIN vccdgt_1p0.gds96
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.446 2.8695 47.502 3.0695 ;
 END
 END vccdgt_1p0.gds96
 PIN vccdgt_1p0.gds97
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.626 3.1075 48.682 3.3075 ;
 END
 END vccdgt_1p0.gds97
 PIN vccdgt_1p0.gds98
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.97 3.1075 50.03 3.3075 ;
 END
 END vccdgt_1p0.gds98
 PIN vccdgt_1p0.gds99
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.606 2.82 47.662 3.02 ;
 END
 END vccdgt_1p0.gds99
 PIN vccdgt_1p0.gds100
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.418 3.1075 49.458 3.3075 ;
 END
 END vccdgt_1p0.gds100
 PIN vccdgt_1p0.gds101
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.266 2.9115 47.342 3.1115 ;
 END
 END vccdgt_1p0.gds101
 PIN vccdgt_1p0.gds102
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.106 3.25 48.182 3.45 ;
 END
 END vccdgt_1p0.gds102
 PIN vccdgt_1p0.gds103
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.29 3.054 49.33 3.254 ;
 END
 END vccdgt_1p0.gds103
 PIN vccdgt_1p0.gds104
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.87 3.054 48.91 3.254 ;
 END
 END vccdgt_1p0.gds104
 PIN vccdgt_1p0.gds105
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.286 3.25 48.342 3.45 ;
 END
 END vccdgt_1p0.gds105
 PIN vccdgt_1p0.gds106
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.626 3.0365 49.686 3.2365 ;
 END
 END vccdgt_1p0.gds106
 PIN vccdgt_1p0.gds107
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.062 3.3775 49.102 3.5775 ;
 END
 END vccdgt_1p0.gds107
 PIN vccdgt_1p0.gds108
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.134 3.265 50.18 3.465 ;
 END
 END vccdgt_1p0.gds108
 PIN vccdgt_1p0.gds109
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.782 3.0175 46.822 3.2175 ;
 END
 END vccdgt_1p0.gds109
 PIN vccdgt_1p0.gds110
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.506 2.9745 46.566 3.1745 ;
 END
 END vccdgt_1p0.gds110
 PIN vccdgt_1p0.gds111
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 48.86 1.013 48.916 1.213 ;
 RECT 50.036 1.076 50.092 1.276 ;
 RECT 50.204 2.273 50.26 2.473 ;
 RECT 48.86 2.273 48.916 2.473 ;
 RECT 48.86 3.533 48.916 3.733 ;
 RECT 50.204 4.793 50.26 4.993 ;
 RECT 48.86 4.793 48.916 4.993 ;
 RECT 48.104 0.896 48.16 1.096 ;
 RECT 48.104 2.156 48.16 2.356 ;
 RECT 48.104 3.416 48.16 3.616 ;
 RECT 48.104 4.676 48.16 4.876 ;
 RECT 49.028 4.36 49.084 4.56 ;
 RECT 49.868 4.436 49.924 4.636 ;
 RECT 49.616 4.688 49.672 4.888 ;
 RECT 50.036 4.856 50.092 5.056 ;
 RECT 49.364 4.775 49.42 4.975 ;
 RECT 48.692 4.793 48.748 4.993 ;
 RECT 48.524 4.78 48.58 4.98 ;
 RECT 49.028 3.1 49.084 3.3 ;
 RECT 49.868 3.176 49.924 3.376 ;
 RECT 49.616 3.428 49.672 3.628 ;
 RECT 50.036 3.596 50.092 3.796 ;
 RECT 50.204 3.533 50.26 3.733 ;
 RECT 48.692 3.533 48.748 3.733 ;
 RECT 48.524 3.52 48.58 3.72 ;
 RECT 49.364 3.515 49.42 3.715 ;
 RECT 49.028 1.84 49.084 2.04 ;
 RECT 49.868 1.916 49.924 2.116 ;
 RECT 49.616 2.168 49.672 2.368 ;
 RECT 50.036 2.336 50.092 2.536 ;
 RECT 49.364 2.255 49.42 2.455 ;
 RECT 48.692 2.273 48.748 2.473 ;
 RECT 48.524 2.26 48.58 2.46 ;
 RECT 49.028 0.58 49.084 0.78 ;
 RECT 49.868 0.656 49.924 0.856 ;
 RECT 49.616 0.908 49.672 1.108 ;
 RECT 49.364 0.995 49.42 1.195 ;
 RECT 48.692 1.013 48.748 1.213 ;
 RECT 50.204 1.013 50.26 1.213 ;
 RECT 48.524 1 48.58 1.2 ;
 END
 END vccdgt_1p0.gds111
 PIN vccdgt_1p0.gds112
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 1.522 50.674 1.722 ;
 END
 END vccdgt_1p0.gds112
 PIN vccdgt_1p0.gds113
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 2.782 50.674 2.982 ;
 END
 END vccdgt_1p0.gds113
 PIN vccdgt_1p0.gds114
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 4.042 50.674 4.242 ;
 END
 END vccdgt_1p0.gds114
 PIN vccdgt_1p0.gds115
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 5.302 50.674 5.502 ;
 END
 END vccdgt_1p0.gds115
 PIN vccdgt_1p0.gds116
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.122 2.862 51.178 3.062 ;
 END
 END vccdgt_1p0.gds116
 PIN vccdgt_1p0.gds117
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.942 2.8695 50.998 3.0695 ;
 END
 END vccdgt_1p0.gds117
 PIN vccdgt_1p0.gds118
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.442 2.8695 51.518 3.0695 ;
 END
 END vccdgt_1p0.gds118
 PIN vccdgt_1p0.gds119
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.778 2.8695 50.838 3.0695 ;
 END
 END vccdgt_1p0.gds119
 PIN vccdgt_1p0.gds120
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.962 3.016 52.002 3.216 ;
 END
 END vccdgt_1p0.gds120
 PIN vccdgt_1p0.gds121
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.702 3.0505 51.758 3.2505 ;
 END
 END vccdgt_1p0.gds121
 PIN vccdgt_1p0.gds122
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.218 2.9745 52.278 3.1745 ;
 END
 END vccdgt_1p0.gds122
 PIN vccdgt_1p0.gds123
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.282 3.016 51.338 3.216 ;
 END
 END vccdgt_1p0.gds123
 PIN vccdgt_1p0.gds124
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.034 2.978 58.074 3.178 ;
 END
 END vccdgt_1p0.gds124
 PIN vccdgt_1p0.gds125
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.762 2.979 57.802 3.179 ;
 END
 END vccdgt_1p0.gds125
 PIN vccdgt_1p0.gds126
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.498 2.8695 64.554 3.0695 ;
 END
 END vccdgt_1p0.gds126
 PIN vccdgt_1p0.gds127
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.658 2.82 64.714 3.02 ;
 END
 END vccdgt_1p0.gds127
 PIN vccdgt_1p0.gds128
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.318 2.9115 64.394 3.1115 ;
 END
 END vccdgt_1p0.gds128
 PIN vccdgt_1p0.gds129
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.158 3.25 65.234 3.45 ;
 END
 END vccdgt_1p0.gds129
 PIN vccdgt_1p0.gds130
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.834 3.0175 63.874 3.2175 ;
 END
 END vccdgt_1p0.gds130
 PIN vccdgt_1p0.gds131
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.558 2.9745 63.618 3.1745 ;
 END
 END vccdgt_1p0.gds131
 PIN vccdgt_1p0.gds132
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 65.156 0.896 65.212 1.096 ;
 RECT 65.156 2.156 65.212 2.356 ;
 RECT 65.156 3.416 65.212 3.616 ;
 RECT 65.156 4.676 65.212 4.876 ;
 END
 END vccdgt_1p0.gds132
 PIN vccdgt_1p0.gds133
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.678 3.1075 65.734 3.3075 ;
 END
 END vccdgt_1p0.gds133
 PIN vccdgt_1p0.gds134
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 1.522 67.726 1.722 ;
 END
 END vccdgt_1p0.gds134
 PIN vccdgt_1p0.gds135
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 2.782 67.726 2.982 ;
 END
 END vccdgt_1p0.gds135
 PIN vccdgt_1p0.gds136
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 4.042 67.726 4.242 ;
 END
 END vccdgt_1p0.gds136
 PIN vccdgt_1p0.gds137
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 5.302 67.726 5.502 ;
 END
 END vccdgt_1p0.gds137
 PIN vccdgt_1p0.gds138
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.174 2.862 68.23 3.062 ;
 END
 END vccdgt_1p0.gds138
 PIN vccdgt_1p0.gds139
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.994 2.8695 68.05 3.0695 ;
 END
 END vccdgt_1p0.gds139
 PIN vccdgt_1p0.gds140
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.022 3.1075 67.082 3.3075 ;
 END
 END vccdgt_1p0.gds140
 PIN vccdgt_1p0.gds141
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.342 3.054 66.382 3.254 ;
 END
 END vccdgt_1p0.gds141
 PIN vccdgt_1p0.gds142
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.922 3.054 65.962 3.254 ;
 END
 END vccdgt_1p0.gds142
 PIN vccdgt_1p0.gds143
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.338 3.25 65.394 3.45 ;
 END
 END vccdgt_1p0.gds143
 PIN vccdgt_1p0.gds144
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.014 3.016 69.054 3.216 ;
 END
 END vccdgt_1p0.gds144
 PIN vccdgt_1p0.gds145
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.678 3.0365 66.738 3.2365 ;
 END
 END vccdgt_1p0.gds145
 PIN vccdgt_1p0.gds146
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.754 3.0505 68.81 3.2505 ;
 END
 END vccdgt_1p0.gds146
 PIN vccdgt_1p0.gds147
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.494 2.8695 68.57 3.0695 ;
 END
 END vccdgt_1p0.gds147
 PIN vccdgt_1p0.gds148
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.83 2.8695 67.89 3.0695 ;
 END
 END vccdgt_1p0.gds148
 PIN vccdgt_1p0.gds149
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.47 3.1075 66.51 3.3075 ;
 END
 END vccdgt_1p0.gds149
 PIN vccdgt_1p0.gds150
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.27 2.9745 69.33 3.1745 ;
 END
 END vccdgt_1p0.gds150
 PIN vccdgt_1p0.gds151
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.334 3.016 68.39 3.216 ;
 END
 END vccdgt_1p0.gds151
 PIN vccdgt_1p0.gds152
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.114 3.3775 66.154 3.5775 ;
 END
 END vccdgt_1p0.gds152
 PIN vccdgt_1p0.gds153
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.186 3.265 67.232 3.465 ;
 END
 END vccdgt_1p0.gds153
 PIN vccdgt_1p0.gds154
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 65.912 1.013 65.968 1.213 ;
 RECT 67.088 1.076 67.144 1.276 ;
 RECT 67.256 2.273 67.312 2.473 ;
 RECT 65.912 2.273 65.968 2.473 ;
 RECT 65.912 3.533 65.968 3.733 ;
 RECT 67.256 4.793 67.312 4.993 ;
 RECT 65.912 4.793 65.968 4.993 ;
 RECT 66.08 4.36 66.136 4.56 ;
 RECT 66.92 4.436 66.976 4.636 ;
 RECT 66.668 4.688 66.724 4.888 ;
 RECT 67.088 4.856 67.144 5.056 ;
 RECT 66.416 4.775 66.472 4.975 ;
 RECT 65.744 4.793 65.8 4.993 ;
 RECT 65.576 4.78 65.632 4.98 ;
 RECT 66.08 3.1 66.136 3.3 ;
 RECT 66.92 3.176 66.976 3.376 ;
 RECT 66.668 3.428 66.724 3.628 ;
 RECT 67.088 3.596 67.144 3.796 ;
 RECT 67.256 3.533 67.312 3.733 ;
 RECT 65.744 3.533 65.8 3.733 ;
 RECT 65.576 3.52 65.632 3.72 ;
 RECT 66.416 3.515 66.472 3.715 ;
 RECT 66.08 1.84 66.136 2.04 ;
 RECT 66.92 1.916 66.976 2.116 ;
 RECT 66.668 2.168 66.724 2.368 ;
 RECT 67.088 2.336 67.144 2.536 ;
 RECT 66.416 2.255 66.472 2.455 ;
 RECT 65.744 2.273 65.8 2.473 ;
 RECT 65.576 2.26 65.632 2.46 ;
 RECT 66.08 0.58 66.136 0.78 ;
 RECT 66.92 0.656 66.976 0.856 ;
 RECT 66.668 0.908 66.724 1.108 ;
 RECT 66.416 0.995 66.472 1.195 ;
 RECT 65.744 1.013 65.8 1.213 ;
 RECT 67.256 1.013 67.312 1.213 ;
 RECT 65.576 1 65.632 1.2 ;
 END
 END vccdgt_1p0.gds154
 PIN vccdgt_1p0.gds155
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 6.239 0.654 6.439 ;
 END
 END vccdgt_1p0.gds155
 PIN vccdgt_1p0.gds156
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 8.759 0.654 8.959 ;
 END
 END vccdgt_1p0.gds156
 PIN vccdgt_1p0.gds157
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 10.019 0.654 10.219 ;
 END
 END vccdgt_1p0.gds157
 PIN vccdgt_1p0.gds158
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 7.499 0.654 7.699 ;
 END
 END vccdgt_1p0.gds158
 PIN vccdgt_1p0.gds159
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.454 8.14 0.494 8.34 ;
 END
 END vccdgt_1p0.gds159
 PIN vccdgt_1p0.gds160
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.742 8.0905 0.788 8.2905 ;
 END
 END vccdgt_1p0.gds160
 PIN vccdgt_1p0.gds161
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.114 8.043 1.154 8.243 ;
 END
 END vccdgt_1p0.gds161
 PIN vccdgt_1p0.gds162
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.566 7.943 1.622 8.143 ;
 END
 END vccdgt_1p0.gds162
 PIN vccdgt_1p0.gds163
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.166 8.006 3.206 8.206 ;
 END
 END vccdgt_1p0.gds163
 PIN vccdgt_1p0.gds164
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.966 8.0065 1.026 8.2065 ;
 END
 END vccdgt_1p0.gds164
 PIN vccdgt_1p0.gds165
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.986 8.0825 2.042 8.2825 ;
 END
 END vccdgt_1p0.gds165
 PIN vccdgt_1p0.gds166
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.326 8.0545 2.382 8.2545 ;
 END
 END vccdgt_1p0.gds166
 PIN vccdgt_1p0.gds167
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.806 8.1355 1.882 8.3355 ;
 END
 END vccdgt_1p0.gds167
 PIN vccdgt_1p0.gds168
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.646 8.0145 2.722 8.2145 ;
 END
 END vccdgt_1p0.gds168
 PIN vccdgt_1p0.gds169
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.634 8.179 4.674 8.379 ;
 END
 END vccdgt_1p0.gds169
 PIN vccdgt_1p0.gds170
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.098 8.0355 5.138 8.2355 ;
 END
 END vccdgt_1p0.gds170
 PIN vccdgt_1p0.gds171
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.478 8.02 3.538 8.22 ;
 END
 END vccdgt_1p0.gds171
 PIN vccdgt_1p0.gds172
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.69 8.099 3.73 8.299 ;
 END
 END vccdgt_1p0.gds172
 PIN vccdgt_1p0.gds173
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.882 8.1125 3.922 8.3125 ;
 END
 END vccdgt_1p0.gds173
 PIN vccdgt_1p0.gds174
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.362 8.165 4.418 8.365 ;
 END
 END vccdgt_1p0.gds174
 PIN vccdgt_1p0.gds175
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.09 8.0905 4.13 8.2905 ;
 END
 END vccdgt_1p0.gds175
 PIN vccdgt_1p0.gds176
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.906 8.122 4.946 8.322 ;
 END
 END vccdgt_1p0.gds176
 PIN vccdgt_1p0.gds177
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.762 8.018 4.818 8.218 ;
 END
 END vccdgt_1p0.gds177
 PIN vccdgt_1p0.gds178
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.486 8.098 2.542 8.298 ;
 END
 END vccdgt_1p0.gds178
 PIN vccdgt_1p0.gds179
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 1.232 6.516 1.288 6.716 ;
 RECT 1.568 6.531 1.624 6.731 ;
 RECT 1.82 6.531 1.876 6.731 ;
 RECT 2.072 6.645 2.128 6.825 ;
 RECT 2.996 6.643 3.052 6.825 ;
 RECT 3.164 6.643 3.22 6.819 ;
 RECT 2.492 6.1445 2.548 6.3445 ;
 RECT 1.232 7.776 1.288 7.976 ;
 RECT 1.568 7.791 1.624 7.991 ;
 RECT 1.82 7.791 1.876 7.991 ;
 RECT 2.072 7.905 2.128 8.085 ;
 RECT 2.996 7.903 3.052 8.085 ;
 RECT 3.164 7.903 3.22 8.079 ;
 RECT 2.492 7.4045 2.548 7.6045 ;
 RECT 1.232 9.036 1.288 9.236 ;
 RECT 1.568 9.051 1.624 9.251 ;
 RECT 1.82 9.051 1.876 9.251 ;
 RECT 2.072 9.165 2.128 9.345 ;
 RECT 2.996 9.163 3.052 9.345 ;
 RECT 3.164 9.163 3.22 9.339 ;
 RECT 2.492 8.6645 2.548 8.8645 ;
 RECT 1.232 10.296 1.288 10.496 ;
 RECT 1.568 10.311 1.624 10.511 ;
 RECT 1.82 10.311 1.876 10.511 ;
 RECT 2.072 10.425 2.128 10.605 ;
 RECT 2.996 10.423 3.052 10.605 ;
 RECT 3.164 10.423 3.22 10.599 ;
 RECT 2.492 9.9245 2.548 10.1245 ;
 RECT 0.812 10.329 0.868 10.529 ;
 RECT 0.644 10.329 0.7 10.529 ;
 RECT 0.98 10.329 1.036 10.529 ;
 RECT 0.812 6.549 0.868 6.749 ;
 RECT 0.644 6.549 0.7 6.749 ;
 RECT 0.98 6.549 1.036 6.749 ;
 RECT 0.812 7.809 0.868 8.009 ;
 RECT 0.644 7.809 0.7 8.009 ;
 RECT 0.98 7.809 1.036 8.009 ;
 RECT 0.812 9.069 0.868 9.269 ;
 RECT 0.644 9.069 0.7 9.269 ;
 RECT 0.98 9.069 1.036 9.269 ;
 RECT 4.088 9.8735 4.144 10.0735 ;
 RECT 4.676 9.8735 4.732 10.0735 ;
 RECT 4.424 9.8735 4.48 10.0735 ;
 RECT 5.012 9.8735 5.068 10.0735 ;
 RECT 4.844 9.8735 4.9 10.0735 ;
 RECT 4.088 8.6135 4.144 8.8135 ;
 RECT 4.676 8.6135 4.732 8.8135 ;
 RECT 4.424 8.6135 4.48 8.8135 ;
 RECT 5.012 8.6135 5.068 8.8135 ;
 RECT 4.844 8.6135 4.9 8.8135 ;
 RECT 4.088 7.3535 4.144 7.5535 ;
 RECT 4.676 7.3535 4.732 7.5535 ;
 RECT 4.424 7.3535 4.48 7.5535 ;
 RECT 5.012 7.3535 5.068 7.5535 ;
 RECT 4.844 7.3535 4.9 7.5535 ;
 RECT 4.088 6.0935 4.144 6.2935 ;
 RECT 4.676 6.0935 4.732 6.2935 ;
 RECT 4.424 6.0935 4.48 6.2935 ;
 RECT 5.012 6.0935 5.068 6.2935 ;
 RECT 4.844 6.0935 4.9 6.2935 ;
 END
 END vccdgt_1p0.gds179
 PIN vccdgt_1p0.gds180
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.33 8.778 6.37 8.978 ;
 END
 END vccdgt_1p0.gds180
 PIN vccdgt_1p0.gds181
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.498 8.02 5.538 8.22 ;
 END
 END vccdgt_1p0.gds181
 PIN vccdgt_1p0.gds182
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.862 8.1125 6.918 8.3125 ;
 END
 END vccdgt_1p0.gds182
 PIN vccdgt_1p0.gds183
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.074 8.122 6.114 8.322 ;
 END
 END vccdgt_1p0.gds183
 PIN vccdgt_1p0.gds184
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.306 8.1125 5.346 8.3125 ;
 END
 END vccdgt_1p0.gds184
 PIN vccdgt_1p0.gds185
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.818 8.0905 5.858 8.2905 ;
 END
 END vccdgt_1p0.gds185
 PIN vccdgt_1p0.gds186
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.626 8.1145 5.666 8.3145 ;
 END
 END vccdgt_1p0.gds186
 PIN vccdgt_1p0.gds187
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.202 8.0995 6.242 8.2995 ;
 END
 END vccdgt_1p0.gds187
 PIN vccdgt_1p0.gds188
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.67 8.039 6.71 8.239 ;
 END
 END vccdgt_1p0.gds188
 PIN vccdgt_1p0.gds189
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.348 9.9245 5.404 10.1245 ;
 RECT 6.02 9.8735 6.076 10.0735 ;
 RECT 5.684 9.9525 5.74 10.1525 ;
 RECT 6.356 9.9525 6.412 10.1525 ;
 RECT 5.348 8.6645 5.404 8.8645 ;
 RECT 6.02 8.6135 6.076 8.8135 ;
 RECT 5.684 8.6925 5.74 8.8925 ;
 RECT 6.356 8.6925 6.412 8.8925 ;
 RECT 5.348 7.4045 5.404 7.6045 ;
 RECT 6.02 7.3535 6.076 7.5535 ;
 RECT 5.684 7.4325 5.74 7.6325 ;
 RECT 6.356 7.4325 6.412 7.6325 ;
 RECT 5.348 6.1445 5.404 6.3445 ;
 RECT 6.02 6.0935 6.076 6.2935 ;
 RECT 5.684 6.1725 5.74 6.3725 ;
 RECT 6.356 6.1725 6.412 6.3725 ;
 END
 END vccdgt_1p0.gds189
 PIN vccdgt_1p0.gds190
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.522 8.8965 14.578 9.0965 ;
 END
 END vccdgt_1p0.gds190
 PIN vccdgt_1p0.gds191
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.342 7.9095 13.398 8.1095 ;
 END
 END vccdgt_1p0.gds191
 PIN vccdgt_1p0.gds192
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.186 8.4265 15.226 8.6265 ;
 END
 END vccdgt_1p0.gds192
 PIN vccdgt_1p0.gds193
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.502 7.86 13.558 8.06 ;
 END
 END vccdgt_1p0.gds193
 PIN vccdgt_1p0.gds194
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.182 8.8105 14.238 9.0105 ;
 END
 END vccdgt_1p0.gds194
 PIN vccdgt_1p0.gds195
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.766 8.094 14.806 8.294 ;
 END
 END vccdgt_1p0.gds195
 PIN vccdgt_1p0.gds196
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.678 8.0575 12.718 8.2575 ;
 END
 END vccdgt_1p0.gds196
 PIN vccdgt_1p0.gds197
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.162 7.9515 13.238 8.1515 ;
 END
 END vccdgt_1p0.gds197
 PIN vccdgt_1p0.gds198
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.002 9.0575 14.078 9.2575 ;
 END
 END vccdgt_1p0.gds198
 PIN vccdgt_1p0.gds199
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.958 9.093 14.998 9.293 ;
 END
 END vccdgt_1p0.gds199
 PIN vccdgt_1p0.gds200
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.402 8.0145 12.462 8.2145 ;
 END
 END vccdgt_1p0.gds200
 PIN vccdgt_1p0.gds201
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 14.756 6.053 14.812 6.253 ;
 RECT 14 7.196 14.056 7.396 ;
 RECT 14.756 7.313 14.812 7.513 ;
 RECT 14 9.716 14.056 9.916 ;
 RECT 14.756 9.833 14.812 10.033 ;
 RECT 14.924 9.4 14.98 9.6 ;
 RECT 14.588 9.833 14.644 10.033 ;
 RECT 14.42 9.82 14.476 10.02 ;
 RECT 14 8.456 14.056 8.656 ;
 RECT 14.756 8.573 14.812 8.773 ;
 RECT 14.924 8.14 14.98 8.34 ;
 RECT 14.588 8.573 14.644 8.773 ;
 RECT 14.42 8.56 14.476 8.76 ;
 RECT 14.924 6.88 14.98 7.08 ;
 RECT 14.588 7.313 14.644 7.513 ;
 RECT 14.42 7.3 14.476 7.5 ;
 RECT 14 5.936 14.056 6.136 ;
 RECT 14.924 5.62 14.98 5.82 ;
 RECT 14.588 6.053 14.644 6.253 ;
 RECT 14.42 6.04 14.476 6.24 ;
 END
 END vccdgt_1p0.gds201
 PIN vccdgt_1p0.gds202
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 6.562 16.57 6.762 ;
 END
 END vccdgt_1p0.gds202
 PIN vccdgt_1p0.gds203
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 7.822 16.57 8.022 ;
 END
 END vccdgt_1p0.gds203
 PIN vccdgt_1p0.gds204
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 9.082 16.57 9.282 ;
 END
 END vccdgt_1p0.gds204
 PIN vccdgt_1p0.gds205
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.018 8.2085 17.074 8.4085 ;
 END
 END vccdgt_1p0.gds205
 PIN vccdgt_1p0.gds206
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.838 7.9095 16.894 8.1095 ;
 END
 END vccdgt_1p0.gds206
 PIN vccdgt_1p0.gds207
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.866 8.8965 15.926 9.0965 ;
 END
 END vccdgt_1p0.gds207
 PIN vccdgt_1p0.gds208
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.03 9.3945 16.076 9.5945 ;
 END
 END vccdgt_1p0.gds208
 PIN vccdgt_1p0.gds209
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.314 8.094 15.354 8.294 ;
 END
 END vccdgt_1p0.gds209
 PIN vccdgt_1p0.gds210
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.338 7.9095 17.414 8.1095 ;
 END
 END vccdgt_1p0.gds210
 PIN vccdgt_1p0.gds211
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.522 8.0765 15.582 8.2765 ;
 END
 END vccdgt_1p0.gds211
 PIN vccdgt_1p0.gds212
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.598 8.0905 17.654 8.2905 ;
 END
 END vccdgt_1p0.gds212
 PIN vccdgt_1p0.gds213
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.674 7.9095 16.734 8.1095 ;
 END
 END vccdgt_1p0.gds213
 PIN vccdgt_1p0.gds214
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.858 8.056 17.898 8.256 ;
 END
 END vccdgt_1p0.gds214
 PIN vccdgt_1p0.gds215
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.114 8.0145 18.174 8.2145 ;
 END
 END vccdgt_1p0.gds215
 PIN vccdgt_1p0.gds216
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.178 8.056 17.234 8.256 ;
 END
 END vccdgt_1p0.gds216
 PIN vccdgt_1p0.gds217
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 16.1 8.573 16.156 8.773 ;
 RECT 15.764 9.476 15.82 9.676 ;
 RECT 15.512 9.728 15.568 9.928 ;
 RECT 15.932 9.896 15.988 10.096 ;
 RECT 16.1 9.833 16.156 10.033 ;
 RECT 15.26 9.815 15.316 10.015 ;
 RECT 15.932 8.636 15.988 8.836 ;
 RECT 15.764 8.216 15.82 8.416 ;
 RECT 15.512 8.468 15.568 8.668 ;
 RECT 15.26 8.555 15.316 8.755 ;
 RECT 15.764 6.956 15.82 7.156 ;
 RECT 15.512 7.208 15.568 7.408 ;
 RECT 15.932 7.376 15.988 7.576 ;
 RECT 16.1 7.313 16.156 7.513 ;
 RECT 15.26 7.295 15.316 7.495 ;
 RECT 15.764 5.696 15.82 5.896 ;
 RECT 15.512 5.948 15.568 6.148 ;
 RECT 15.932 6.116 15.988 6.316 ;
 RECT 16.1 6.053 16.156 6.253 ;
 RECT 15.26 6.035 15.316 6.235 ;
 END
 END vccdgt_1p0.gds217
 PIN vccdgt_1p0.gds218
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.93 8.018 23.97 8.218 ;
 END
 END vccdgt_1p0.gds218
 PIN vccdgt_1p0.gds219
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.658 8.019 23.698 8.219 ;
 END
 END vccdgt_1p0.gds219
 PIN vccdgt_1p0.gds220
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.214 7.9515 30.29 8.1515 ;
 END
 END vccdgt_1p0.gds220
 PIN vccdgt_1p0.gds221
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.73 8.0575 29.77 8.2575 ;
 END
 END vccdgt_1p0.gds221
 PIN vccdgt_1p0.gds222
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.454 8.0145 29.514 8.2145 ;
 END
 END vccdgt_1p0.gds222
 PIN vccdgt_1p0.gds223
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 7.822 33.622 8.022 ;
 END
 END vccdgt_1p0.gds223
 PIN vccdgt_1p0.gds224
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 6.562 33.622 6.762 ;
 END
 END vccdgt_1p0.gds224
 PIN vccdgt_1p0.gds225
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 9.082 33.622 9.282 ;
 END
 END vccdgt_1p0.gds225
 PIN vccdgt_1p0.gds226
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.07 8.2085 34.126 8.4085 ;
 END
 END vccdgt_1p0.gds226
 PIN vccdgt_1p0.gds227
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.89 7.9095 33.946 8.1095 ;
 END
 END vccdgt_1p0.gds227
 PIN vccdgt_1p0.gds228
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.918 8.8965 32.978 9.0965 ;
 END
 END vccdgt_1p0.gds228
 PIN vccdgt_1p0.gds229
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.574 8.8965 31.63 9.0965 ;
 END
 END vccdgt_1p0.gds229
 PIN vccdgt_1p0.gds230
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.394 7.9095 30.45 8.1095 ;
 END
 END vccdgt_1p0.gds230
 PIN vccdgt_1p0.gds231
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.39 7.9095 34.466 8.1095 ;
 END
 END vccdgt_1p0.gds231
 PIN vccdgt_1p0.gds232
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.238 8.094 32.278 8.294 ;
 END
 END vccdgt_1p0.gds232
 PIN vccdgt_1p0.gds233
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.818 8.094 31.858 8.294 ;
 END
 END vccdgt_1p0.gds233
 PIN vccdgt_1p0.gds234
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.234 8.8105 31.29 9.0105 ;
 END
 END vccdgt_1p0.gds234
 PIN vccdgt_1p0.gds235
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.082 9.3945 33.128 9.5945 ;
 END
 END vccdgt_1p0.gds235
 PIN vccdgt_1p0.gds236
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.366 8.4265 32.406 8.6265 ;
 END
 END vccdgt_1p0.gds236
 PIN vccdgt_1p0.gds237
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.01 9.093 32.05 9.293 ;
 END
 END vccdgt_1p0.gds237
 PIN vccdgt_1p0.gds238
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.166 8.0145 35.226 8.2145 ;
 END
 END vccdgt_1p0.gds238
 PIN vccdgt_1p0.gds239
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.91 8.056 34.95 8.256 ;
 END
 END vccdgt_1p0.gds239
 PIN vccdgt_1p0.gds240
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.054 9.0575 31.13 9.2575 ;
 END
 END vccdgt_1p0.gds240
 PIN vccdgt_1p0.gds241
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.554 7.86 30.61 8.06 ;
 END
 END vccdgt_1p0.gds241
 PIN vccdgt_1p0.gds242
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.23 8.056 34.286 8.256 ;
 END
 END vccdgt_1p0.gds242
 PIN vccdgt_1p0.gds243
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.65 8.0905 34.706 8.2905 ;
 END
 END vccdgt_1p0.gds243
 PIN vccdgt_1p0.gds244
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.574 8.0765 32.634 8.2765 ;
 END
 END vccdgt_1p0.gds244
 PIN vccdgt_1p0.gds245
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.726 7.9095 33.786 8.1095 ;
 END
 END vccdgt_1p0.gds245
 PIN vccdgt_1p0.gds246
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 33.152 6.053 33.208 6.253 ;
 RECT 31.808 9.833 31.864 10.033 ;
 RECT 32.984 9.896 33.04 10.096 ;
 RECT 31.976 9.4 32.032 9.6 ;
 RECT 32.816 9.476 32.872 9.676 ;
 RECT 33.152 8.573 33.208 8.773 ;
 RECT 33.152 7.313 33.208 7.513 ;
 RECT 31.808 7.313 31.864 7.513 ;
 RECT 31.808 8.573 31.864 8.773 ;
 RECT 31.052 7.196 31.108 7.396 ;
 RECT 31.052 8.456 31.108 8.656 ;
 RECT 31.052 9.716 31.108 9.916 ;
 RECT 31.976 8.14 32.032 8.34 ;
 RECT 32.816 8.216 32.872 8.416 ;
 RECT 32.564 8.468 32.62 8.668 ;
 RECT 32.984 8.636 33.04 8.836 ;
 RECT 31.976 6.88 32.032 7.08 ;
 RECT 32.816 6.956 32.872 7.156 ;
 RECT 32.564 7.208 32.62 7.408 ;
 RECT 32.984 7.376 33.04 7.576 ;
 RECT 32.312 7.295 32.368 7.495 ;
 RECT 31.64 7.313 31.696 7.513 ;
 RECT 31.472 7.3 31.528 7.5 ;
 RECT 32.312 8.555 32.368 8.755 ;
 RECT 31.64 8.573 31.696 8.773 ;
 RECT 31.472 8.56 31.528 8.76 ;
 RECT 32.564 9.728 32.62 9.928 ;
 RECT 32.312 9.815 32.368 10.015 ;
 RECT 31.64 9.833 31.696 10.033 ;
 RECT 33.152 9.833 33.208 10.033 ;
 RECT 31.472 9.82 31.528 10.02 ;
 RECT 31.052 5.936 31.108 6.136 ;
 RECT 31.808 6.053 31.864 6.253 ;
 RECT 32.984 6.116 33.04 6.316 ;
 RECT 31.976 5.62 32.032 5.82 ;
 RECT 32.816 5.696 32.872 5.896 ;
 RECT 32.564 5.948 32.62 6.148 ;
 RECT 32.312 6.035 32.368 6.235 ;
 RECT 31.64 6.053 31.696 6.253 ;
 RECT 31.472 6.04 31.528 6.24 ;
 END
 END vccdgt_1p0.gds246
 PIN vccdgt_1p0.gds247
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.982 8.018 41.022 8.218 ;
 END
 END vccdgt_1p0.gds247
 PIN vccdgt_1p0.gds248
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.71 8.019 40.75 8.219 ;
 END
 END vccdgt_1p0.gds248
 PIN vccdgt_1p0.gds249
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.446 7.9095 47.502 8.1095 ;
 END
 END vccdgt_1p0.gds249
 PIN vccdgt_1p0.gds250
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.626 8.8965 48.682 9.0965 ;
 END
 END vccdgt_1p0.gds250
 PIN vccdgt_1p0.gds251
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.97 8.8965 50.03 9.0965 ;
 END
 END vccdgt_1p0.gds251
 PIN vccdgt_1p0.gds252
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.606 7.86 47.662 8.06 ;
 END
 END vccdgt_1p0.gds252
 PIN vccdgt_1p0.gds253
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.418 8.4265 49.458 8.6265 ;
 END
 END vccdgt_1p0.gds253
 PIN vccdgt_1p0.gds254
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.266 7.9515 47.342 8.1515 ;
 END
 END vccdgt_1p0.gds254
 PIN vccdgt_1p0.gds255
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.106 9.0575 48.182 9.2575 ;
 END
 END vccdgt_1p0.gds255
 PIN vccdgt_1p0.gds256
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.29 8.094 49.33 8.294 ;
 END
 END vccdgt_1p0.gds256
 PIN vccdgt_1p0.gds257
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.87 8.094 48.91 8.294 ;
 END
 END vccdgt_1p0.gds257
 PIN vccdgt_1p0.gds258
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.286 8.8105 48.342 9.0105 ;
 END
 END vccdgt_1p0.gds258
 PIN vccdgt_1p0.gds259
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.626 8.0765 49.686 8.2765 ;
 END
 END vccdgt_1p0.gds259
 PIN vccdgt_1p0.gds260
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.062 9.093 49.102 9.293 ;
 END
 END vccdgt_1p0.gds260
 PIN vccdgt_1p0.gds261
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.134 9.3945 50.18 9.5945 ;
 END
 END vccdgt_1p0.gds261
 PIN vccdgt_1p0.gds262
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.782 8.0575 46.822 8.2575 ;
 END
 END vccdgt_1p0.gds262
 PIN vccdgt_1p0.gds263
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.506 8.0145 46.566 8.2145 ;
 END
 END vccdgt_1p0.gds263
 PIN vccdgt_1p0.gds264
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 50.204 6.053 50.26 6.253 ;
 RECT 48.104 7.196 48.16 7.396 ;
 RECT 48.86 7.313 48.916 7.513 ;
 RECT 50.204 8.573 50.26 8.773 ;
 RECT 48.104 9.716 48.16 9.916 ;
 RECT 48.86 9.833 48.916 10.033 ;
 RECT 49.028 9.4 49.084 9.6 ;
 RECT 49.868 9.476 49.924 9.676 ;
 RECT 49.616 9.728 49.672 9.928 ;
 RECT 50.036 9.896 50.092 10.096 ;
 RECT 48.692 9.833 48.748 10.033 ;
 RECT 50.204 9.833 50.26 10.033 ;
 RECT 48.524 9.82 48.58 10.02 ;
 RECT 49.364 9.815 49.42 10.015 ;
 RECT 48.104 8.456 48.16 8.656 ;
 RECT 48.86 8.573 48.916 8.773 ;
 RECT 50.036 8.636 50.092 8.836 ;
 RECT 49.028 8.14 49.084 8.34 ;
 RECT 49.868 8.216 49.924 8.416 ;
 RECT 49.616 8.468 49.672 8.668 ;
 RECT 49.364 8.555 49.42 8.755 ;
 RECT 48.692 8.573 48.748 8.773 ;
 RECT 48.524 8.56 48.58 8.76 ;
 RECT 49.028 6.88 49.084 7.08 ;
 RECT 49.868 6.956 49.924 7.156 ;
 RECT 49.616 7.208 49.672 7.408 ;
 RECT 50.036 7.376 50.092 7.576 ;
 RECT 48.692 7.313 48.748 7.513 ;
 RECT 50.204 7.313 50.26 7.513 ;
 RECT 48.524 7.3 48.58 7.5 ;
 RECT 49.364 7.295 49.42 7.495 ;
 RECT 48.104 5.936 48.16 6.136 ;
 RECT 48.86 6.053 48.916 6.253 ;
 RECT 50.036 6.116 50.092 6.316 ;
 RECT 49.028 5.62 49.084 5.82 ;
 RECT 49.868 5.696 49.924 5.896 ;
 RECT 49.616 5.948 49.672 6.148 ;
 RECT 49.364 6.035 49.42 6.235 ;
 RECT 48.692 6.053 48.748 6.253 ;
 RECT 48.524 6.04 48.58 6.24 ;
 END
 END vccdgt_1p0.gds264
 PIN vccdgt_1p0.gds265
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 6.562 50.674 6.762 ;
 END
 END vccdgt_1p0.gds265
 PIN vccdgt_1p0.gds266
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 7.822 50.674 8.022 ;
 END
 END vccdgt_1p0.gds266
 PIN vccdgt_1p0.gds267
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 9.082 50.674 9.282 ;
 END
 END vccdgt_1p0.gds267
 PIN vccdgt_1p0.gds268
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.122 8.2085 51.178 8.4085 ;
 END
 END vccdgt_1p0.gds268
 PIN vccdgt_1p0.gds269
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.942 7.9095 50.998 8.1095 ;
 END
 END vccdgt_1p0.gds269
 PIN vccdgt_1p0.gds270
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.442 7.9095 51.518 8.1095 ;
 END
 END vccdgt_1p0.gds270
 PIN vccdgt_1p0.gds271
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.778 7.9095 50.838 8.1095 ;
 END
 END vccdgt_1p0.gds271
 PIN vccdgt_1p0.gds272
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.962 8.056 52.002 8.256 ;
 END
 END vccdgt_1p0.gds272
 PIN vccdgt_1p0.gds273
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.702 8.0905 51.758 8.2905 ;
 END
 END vccdgt_1p0.gds273
 PIN vccdgt_1p0.gds274
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.218 8.0145 52.278 8.2145 ;
 END
 END vccdgt_1p0.gds274
 PIN vccdgt_1p0.gds275
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.282 8.056 51.338 8.256 ;
 END
 END vccdgt_1p0.gds275
 PIN vccdgt_1p0.gds276
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.034 8.018 58.074 8.218 ;
 END
 END vccdgt_1p0.gds276
 PIN vccdgt_1p0.gds277
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.762 8.019 57.802 8.219 ;
 END
 END vccdgt_1p0.gds277
 PIN vccdgt_1p0.gds278
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.498 7.9095 64.554 8.1095 ;
 END
 END vccdgt_1p0.gds278
 PIN vccdgt_1p0.gds279
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.658 7.86 64.714 8.06 ;
 END
 END vccdgt_1p0.gds279
 PIN vccdgt_1p0.gds280
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.318 7.9515 64.394 8.1515 ;
 END
 END vccdgt_1p0.gds280
 PIN vccdgt_1p0.gds281
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.158 9.0575 65.234 9.2575 ;
 END
 END vccdgt_1p0.gds281
 PIN vccdgt_1p0.gds282
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.834 8.0575 63.874 8.2575 ;
 END
 END vccdgt_1p0.gds282
 PIN vccdgt_1p0.gds283
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.558 8.0145 63.618 8.2145 ;
 END
 END vccdgt_1p0.gds283
 PIN vccdgt_1p0.gds284
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 65.156 7.196 65.212 7.396 ;
 RECT 65.156 9.716 65.212 9.916 ;
 RECT 65.156 8.456 65.212 8.656 ;
 RECT 65.156 5.936 65.212 6.136 ;
 END
 END vccdgt_1p0.gds284
 PIN vccdgt_1p0.gds285
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.678 8.8965 65.734 9.0965 ;
 END
 END vccdgt_1p0.gds285
 PIN vccdgt_1p0.gds286
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 6.562 67.726 6.762 ;
 END
 END vccdgt_1p0.gds286
 PIN vccdgt_1p0.gds287
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 7.822 67.726 8.022 ;
 END
 END vccdgt_1p0.gds287
 PIN vccdgt_1p0.gds288
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 9.082 67.726 9.282 ;
 END
 END vccdgt_1p0.gds288
 PIN vccdgt_1p0.gds289
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.174 8.2085 68.23 8.4085 ;
 END
 END vccdgt_1p0.gds289
 PIN vccdgt_1p0.gds290
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.994 7.9095 68.05 8.1095 ;
 END
 END vccdgt_1p0.gds290
 PIN vccdgt_1p0.gds291
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.022 8.8965 67.082 9.0965 ;
 END
 END vccdgt_1p0.gds291
 PIN vccdgt_1p0.gds292
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.342 8.094 66.382 8.294 ;
 END
 END vccdgt_1p0.gds292
 PIN vccdgt_1p0.gds293
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.922 8.094 65.962 8.294 ;
 END
 END vccdgt_1p0.gds293
 PIN vccdgt_1p0.gds294
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.338 8.8105 65.394 9.0105 ;
 END
 END vccdgt_1p0.gds294
 PIN vccdgt_1p0.gds295
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.014 8.056 69.054 8.256 ;
 END
 END vccdgt_1p0.gds295
 PIN vccdgt_1p0.gds296
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.678 8.0765 66.738 8.2765 ;
 END
 END vccdgt_1p0.gds296
 PIN vccdgt_1p0.gds297
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.754 8.0905 68.81 8.2905 ;
 END
 END vccdgt_1p0.gds297
 PIN vccdgt_1p0.gds298
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.494 7.9095 68.57 8.1095 ;
 END
 END vccdgt_1p0.gds298
 PIN vccdgt_1p0.gds299
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.83 7.9095 67.89 8.1095 ;
 END
 END vccdgt_1p0.gds299
 PIN vccdgt_1p0.gds300
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.47 8.4265 66.51 8.6265 ;
 END
 END vccdgt_1p0.gds300
 PIN vccdgt_1p0.gds301
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.27 8.0145 69.33 8.2145 ;
 END
 END vccdgt_1p0.gds301
 PIN vccdgt_1p0.gds302
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.334 8.056 68.39 8.256 ;
 END
 END vccdgt_1p0.gds302
 PIN vccdgt_1p0.gds303
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.114 9.093 66.154 9.293 ;
 END
 END vccdgt_1p0.gds303
 PIN vccdgt_1p0.gds304
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.186 9.3945 67.232 9.5945 ;
 END
 END vccdgt_1p0.gds304
 PIN vccdgt_1p0.gds305
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 67.256 6.053 67.312 6.253 ;
 RECT 65.912 7.313 65.968 7.513 ;
 RECT 67.256 8.573 67.312 8.773 ;
 RECT 65.912 9.833 65.968 10.033 ;
 RECT 66.08 9.4 66.136 9.6 ;
 RECT 66.92 9.476 66.976 9.676 ;
 RECT 66.668 9.728 66.724 9.928 ;
 RECT 67.088 9.896 67.144 10.096 ;
 RECT 65.744 9.833 65.8 10.033 ;
 RECT 67.256 9.833 67.312 10.033 ;
 RECT 65.576 9.82 65.632 10.02 ;
 RECT 66.416 9.815 66.472 10.015 ;
 RECT 65.912 8.573 65.968 8.773 ;
 RECT 67.088 8.636 67.144 8.836 ;
 RECT 66.08 8.14 66.136 8.34 ;
 RECT 66.92 8.216 66.976 8.416 ;
 RECT 66.668 8.468 66.724 8.668 ;
 RECT 66.416 8.555 66.472 8.755 ;
 RECT 65.744 8.573 65.8 8.773 ;
 RECT 65.576 8.56 65.632 8.76 ;
 RECT 66.08 6.88 66.136 7.08 ;
 RECT 66.92 6.956 66.976 7.156 ;
 RECT 66.668 7.208 66.724 7.408 ;
 RECT 67.088 7.376 67.144 7.576 ;
 RECT 65.744 7.313 65.8 7.513 ;
 RECT 67.256 7.313 67.312 7.513 ;
 RECT 65.576 7.3 65.632 7.5 ;
 RECT 66.416 7.295 66.472 7.495 ;
 RECT 65.912 6.053 65.968 6.253 ;
 RECT 67.088 6.116 67.144 6.316 ;
 RECT 66.08 5.62 66.136 5.82 ;
 RECT 66.92 5.696 66.976 5.896 ;
 RECT 66.668 5.948 66.724 6.148 ;
 RECT 66.416 6.035 66.472 6.235 ;
 RECT 65.744 6.053 65.8 6.253 ;
 RECT 65.576 6.04 65.632 6.24 ;
 END
 END vccdgt_1p0.gds305
 PIN vccdgt_1p0.gds306
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 12.393 2.202 12.593 ;
 END
 END vccdgt_1p0.gds306
 PIN vccdgt_1p0.gds307
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 13.669 0.654 13.869 ;
 END
 END vccdgt_1p0.gds307
 PIN vccdgt_1p0.gds308
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.454 13.2555 0.494 13.4555 ;
 END
 END vccdgt_1p0.gds308
 PIN vccdgt_1p0.gds309
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.742 13.118 0.788 13.318 ;
 END
 END vccdgt_1p0.gds309
 PIN vccdgt_1p0.gds310
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.114 13.1015 1.154 13.3015 ;
 END
 END vccdgt_1p0.gds310
 PIN vccdgt_1p0.gds311
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.566 12.8615 1.622 13.0615 ;
 END
 END vccdgt_1p0.gds311
 PIN vccdgt_1p0.gds312
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.166 11.006 3.206 11.206 ;
 END
 END vccdgt_1p0.gds312
 PIN vccdgt_1p0.gds313
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.966 13.227 1.026 13.427 ;
 END
 END vccdgt_1p0.gds313
 PIN vccdgt_1p0.gds314
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.986 13.9275 2.042 14.1275 ;
 END
 END vccdgt_1p0.gds314
 PIN vccdgt_1p0.gds315
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.326 13.03 2.382 13.23 ;
 END
 END vccdgt_1p0.gds315
 PIN vccdgt_1p0.gds316
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.806 13.1325 1.882 13.3325 ;
 END
 END vccdgt_1p0.gds316
 PIN vccdgt_1p0.gds317
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.646 13.243 2.722 13.443 ;
 END
 END vccdgt_1p0.gds317
 PIN vccdgt_1p0.gds318
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.098 15.1185 5.138 15.3185 ;
 END
 END vccdgt_1p0.gds318
 PIN vccdgt_1p0.gds319
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.634 12.868 4.674 13.068 ;
 END
 END vccdgt_1p0.gds319
 PIN vccdgt_1p0.gds320
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.478 13.2855 3.538 13.4855 ;
 END
 END vccdgt_1p0.gds320
 PIN vccdgt_1p0.gds321
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.69 13.1145 3.73 13.3145 ;
 END
 END vccdgt_1p0.gds321
 PIN vccdgt_1p0.gds322
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.882 10.697 3.922 10.897 ;
 END
 END vccdgt_1p0.gds322
 PIN vccdgt_1p0.gds323
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.362 13.3475 4.418 13.5475 ;
 END
 END vccdgt_1p0.gds323
 PIN vccdgt_1p0.gds324
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.09 11.5505 4.13 11.7505 ;
 END
 END vccdgt_1p0.gds324
 PIN vccdgt_1p0.gds325
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.906 10.477 4.946 10.677 ;
 END
 END vccdgt_1p0.gds325
 PIN vccdgt_1p0.gds326
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.762 12.653 4.818 12.853 ;
 END
 END vccdgt_1p0.gds326
 PIN vccdgt_1p0.gds327
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.486 13.1795 2.542 13.3795 ;
 END
 END vccdgt_1p0.gds327
 PIN vccdgt_1p0.gds328
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 3.248 15.129 3.304 15.293 ;
 RECT 4.004 15.129 4.06 15.293 ;
 RECT 3.752 15.129 3.808 15.293 ;
 RECT 0.896 15.09 0.952 15.29 ;
 RECT 0.56 15.09 0.616 15.29 ;
 RECT 1.568 15.09 1.624 15.29 ;
 RECT 1.4 15.09 1.456 15.29 ;
 RECT 2.828 15.09 2.884 15.29 ;
 RECT 2.66 15.09 2.716 15.29 ;
 RECT 4.256 15.127 4.312 15.309 ;
 RECT 4.928 15.127 4.984 15.309 ;
 RECT 3.668 15.351 3.724 15.533 ;
 RECT 3.248 15.369 3.304 15.569 ;
 RECT 3.5 15.2285 3.556 15.4285 ;
 RECT 4.088 15.37 4.144 15.57 ;
 RECT 3.92 15.37 3.976 15.57 ;
 RECT 0.896 15.37 0.952 15.57 ;
 RECT 0.56 15.37 0.616 15.57 ;
 RECT 1.568 15.37 1.624 15.57 ;
 RECT 1.4 15.37 1.456 15.57 ;
 RECT 1.82 15.35 1.876 15.533 ;
 RECT 3.08 15.37 3.136 15.57 ;
 RECT 3.164 13.747 3.22 13.947 ;
 RECT 0.896 13.746 0.952 13.946 ;
 RECT 0.56 13.746 0.616 13.946 ;
 RECT 1.568 13.746 1.624 13.946 ;
 RECT 1.4 13.746 1.456 13.946 ;
 RECT 2.576 13.746 2.632 13.946 ;
 RECT 2.156 13.746 2.212 13.946 ;
 RECT 1.988 13.783 2.044 13.965 ;
 RECT 2.324 13.783 2.38 13.965 ;
 RECT 2.912 13.746 2.968 13.946 ;
 RECT 2.744 13.746 2.8 13.946 ;
 RECT 4.928 13.783 4.984 13.965 ;
 RECT 3.164 12.681 3.22 12.881 ;
 RECT 4.004 11.338 4.06 11.538 ;
 RECT 4.508 11.335 4.564 11.499 ;
 RECT 0.896 11.338 0.952 11.538 ;
 RECT 0.56 11.338 0.616 11.538 ;
 RECT 1.568 11.338 1.624 11.538 ;
 RECT 1.4 11.338 1.456 11.538 ;
 RECT 2.156 11.338 2.212 11.538 ;
 RECT 4.424 11.058 4.48 11.258 ;
 RECT 4.256 11.1965 4.312 11.3965 ;
 RECT 4.76 11.1965 4.816 11.3965 ;
 RECT 5.18 11.1965 5.236 11.3965 ;
 RECT 4.928 11.198 4.984 11.398 ;
 RECT 3.836 11.095 3.892 11.277 ;
 RECT 3.584 11.198 3.64 11.398 ;
 RECT 3.416 11.058 3.472 11.258 ;
 RECT 4.004 11.058 4.06 11.258 ;
 RECT 2.408 11.059 2.464 11.259 ;
 RECT 2.912 11.059 2.968 11.259 ;
 RECT 2.156 11.059 2.212 11.259 ;
 RECT 2.66 11.059 2.716 11.259 ;
 RECT 1.904 11.059 1.96 11.259 ;
 RECT 1.568 11.058 1.624 11.258 ;
 RECT 1.4 11.058 1.456 11.258 ;
 RECT 0.896 11.058 0.952 11.258 ;
 RECT 0.56 11.058 0.616 11.258 ;
 RECT 3.164 11.198 3.22 11.398 ;
 RECT 2.66 11.338 2.716 11.538 ;
 RECT 3.164 12.403 3.22 12.603 ;
 RECT 3.584 12.5405 3.64 12.7405 ;
 RECT 3.416 12.5405 3.472 12.7405 ;
 RECT 4.004 12.542 4.06 12.742 ;
 RECT 3.836 12.542 3.892 12.742 ;
 RECT 4.508 12.5405 4.564 12.7405 ;
 RECT 4.256 12.5405 4.312 12.7405 ;
 RECT 4.76 12.5405 4.816 12.7405 ;
 RECT 5.18 12.5405 5.236 12.7405 ;
 RECT 4.928 12.542 4.984 12.742 ;
 RECT 0.896 12.402 0.952 12.602 ;
 RECT 0.56 12.402 0.616 12.602 ;
 RECT 1.568 12.402 1.624 12.602 ;
 RECT 1.4 12.402 1.456 12.602 ;
 RECT 2.156 12.402 2.212 12.602 ;
 RECT 2.66 12.402 2.716 12.602 ;
 RECT 0.896 12.682 0.952 12.882 ;
 RECT 0.56 12.682 0.616 12.882 ;
 RECT 1.568 12.682 1.624 12.882 ;
 RECT 1.4 12.682 1.456 12.882 ;
 RECT 2.24 12.682 2.296 12.882 ;
 RECT 2.744 12.681 2.8 12.881 ;
 RECT 3.164 14.025 3.22 14.225 ;
 RECT 3.584 13.8845 3.64 14.0845 ;
 RECT 3.416 13.8845 3.472 14.0845 ;
 RECT 4.004 13.886 4.06 14.086 ;
 RECT 3.836 13.886 3.892 14.086 ;
 RECT 0.896 14.026 0.952 14.226 ;
 RECT 0.56 14.026 0.616 14.226 ;
 RECT 1.568 14.026 1.624 14.226 ;
 RECT 1.4 14.026 1.456 14.226 ;
 RECT 2.156 14.026 2.212 14.226 ;
 RECT 1.988 14.026 2.044 14.226 ;
 RECT 1.82 14.026 1.876 14.226 ;
 RECT 2.492 14.026 2.548 14.226 ;
 RECT 2.324 14.026 2.38 14.226 ;
 RECT 5.18 13.886 5.236 14.086 ;
 RECT 4.256 13.8845 4.312 14.0845 ;
 RECT 4.424 13.8845 4.48 14.0845 ;
 RECT 4.928 14.007 4.984 14.189 ;
 RECT 4.676 13.886 4.732 14.086 ;
 RECT 2.156 15.323 2.212 15.523 ;
 RECT 1.988 15.44 2.044 15.64 ;
 RECT 2.492 15.323 2.548 15.523 ;
 RECT 2.324 15.323 2.38 15.523 ;
 RECT 2.912 15.44 2.968 15.64 ;
 RECT 2.744 15.44 2.8 15.64 ;
 RECT 5.18 15.23 5.236 15.43 ;
 RECT 4.424 15.2285 4.48 15.4285 ;
 RECT 4.928 15.351 4.984 15.533 ;
 RECT 4.676 15.23 4.732 15.43 ;
 END
 END vccdgt_1p0.gds328
 PIN vccdgt_1p0.gds329
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.966 11.011 10.026 11.211 ;
 END
 END vccdgt_1p0.gds329
 PIN vccdgt_1p0.gds330
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.798 11.011 9.858 11.211 ;
 END
 END vccdgt_1p0.gds330
 PIN vccdgt_1p0.gds331
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.134 11.011 10.194 11.211 ;
 END
 END vccdgt_1p0.gds331
 PIN vccdgt_1p0.gds332
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.294 11.011 9.354 11.211 ;
 END
 END vccdgt_1p0.gds332
 PIN vccdgt_1p0.gds333
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.126 11.011 9.186 11.211 ;
 END
 END vccdgt_1p0.gds333
 PIN vccdgt_1p0.gds334
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.462 11.011 9.522 11.211 ;
 END
 END vccdgt_1p0.gds334
 PIN vccdgt_1p0.gds335
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.622 11.011 8.682 11.211 ;
 END
 END vccdgt_1p0.gds335
 PIN vccdgt_1p0.gds336
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.454 11.011 8.514 11.211 ;
 END
 END vccdgt_1p0.gds336
 PIN vccdgt_1p0.gds337
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.79 11.011 8.85 11.211 ;
 END
 END vccdgt_1p0.gds337
 PIN vccdgt_1p0.gds338
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.95 11.011 8.01 11.211 ;
 END
 END vccdgt_1p0.gds338
 PIN vccdgt_1p0.gds339
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.782 11.011 7.842 11.211 ;
 END
 END vccdgt_1p0.gds339
 PIN vccdgt_1p0.gds340
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.118 11.011 8.178 11.211 ;
 END
 END vccdgt_1p0.gds340
 PIN vccdgt_1p0.gds341
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.11 11.011 7.17 11.211 ;
 END
 END vccdgt_1p0.gds341
 PIN vccdgt_1p0.gds342
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.278 11.011 7.338 11.211 ;
 END
 END vccdgt_1p0.gds342
 PIN vccdgt_1p0.gds343
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.446 11.011 7.506 11.211 ;
 END
 END vccdgt_1p0.gds343
 PIN vccdgt_1p0.gds344
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.714 12.7505 9.754 12.9505 ;
 END
 END vccdgt_1p0.gds344
 PIN vccdgt_1p0.gds345
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.042 12.7505 9.082 12.9505 ;
 END
 END vccdgt_1p0.gds345
 PIN vccdgt_1p0.gds346
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.37 12.7505 8.41 12.9505 ;
 END
 END vccdgt_1p0.gds346
 PIN vccdgt_1p0.gds347
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.698 12.7505 7.738 12.9505 ;
 END
 END vccdgt_1p0.gds347
 PIN vccdgt_1p0.gds348
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.026 12.7505 7.066 12.9505 ;
 END
 END vccdgt_1p0.gds348
 PIN vccdgt_1p0.gds349
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.33 13.4825 6.37 13.6825 ;
 END
 END vccdgt_1p0.gds349
 PIN vccdgt_1p0.gds350
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.11 11.9905 10.15 12.1905 ;
 END
 END vccdgt_1p0.gds350
 PIN vccdgt_1p0.gds351
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.438 11.9905 9.478 12.1905 ;
 END
 END vccdgt_1p0.gds351
 PIN vccdgt_1p0.gds352
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.766 11.9905 8.806 12.1905 ;
 END
 END vccdgt_1p0.gds352
 PIN vccdgt_1p0.gds353
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.094 11.9905 8.134 12.1905 ;
 END
 END vccdgt_1p0.gds353
 PIN vccdgt_1p0.gds354
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.498 11.695 5.538 11.895 ;
 END
 END vccdgt_1p0.gds354
 PIN vccdgt_1p0.gds355
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.11 15.406 10.15 15.606 ;
 END
 END vccdgt_1p0.gds355
 PIN vccdgt_1p0.gds356
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.438 15.406 9.478 15.606 ;
 END
 END vccdgt_1p0.gds356
 PIN vccdgt_1p0.gds357
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.766 15.406 8.806 15.606 ;
 END
 END vccdgt_1p0.gds357
 PIN vccdgt_1p0.gds358
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.094 15.406 8.134 15.606 ;
 END
 END vccdgt_1p0.gds358
 PIN vccdgt_1p0.gds359
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.422 15.406 7.462 15.606 ;
 END
 END vccdgt_1p0.gds359
 PIN vccdgt_1p0.gds360
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.918 12.617 9.958 12.817 ;
 END
 END vccdgt_1p0.gds360
 PIN vccdgt_1p0.gds361
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.566 13.483 9.606 13.683 ;
 END
 END vccdgt_1p0.gds361
 PIN vccdgt_1p0.gds362
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.894 13.483 8.934 13.683 ;
 END
 END vccdgt_1p0.gds362
 PIN vccdgt_1p0.gds363
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.246 12.617 9.286 12.817 ;
 END
 END vccdgt_1p0.gds363
 PIN vccdgt_1p0.gds364
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.222 13.483 8.262 13.683 ;
 END
 END vccdgt_1p0.gds364
 PIN vccdgt_1p0.gds365
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.574 12.617 8.614 12.817 ;
 END
 END vccdgt_1p0.gds365
 PIN vccdgt_1p0.gds366
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.23 12.617 7.27 12.817 ;
 END
 END vccdgt_1p0.gds366
 PIN vccdgt_1p0.gds367
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.902 12.617 7.942 12.817 ;
 END
 END vccdgt_1p0.gds367
 PIN vccdgt_1p0.gds368
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.55 13.483 7.59 13.683 ;
 END
 END vccdgt_1p0.gds368
 PIN vccdgt_1p0.gds369
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.862 13.1165 6.918 13.3165 ;
 END
 END vccdgt_1p0.gds369
 PIN vccdgt_1p0.gds370
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.074 13.0285 6.114 13.2285 ;
 END
 END vccdgt_1p0.gds370
 PIN vccdgt_1p0.gds371
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.306 13.1805 5.346 13.3805 ;
 END
 END vccdgt_1p0.gds371
 PIN vccdgt_1p0.gds372
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.818 12.793 5.858 12.993 ;
 END
 END vccdgt_1p0.gds372
 PIN vccdgt_1p0.gds373
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.626 11.1105 5.666 11.3105 ;
 END
 END vccdgt_1p0.gds373
 PIN vccdgt_1p0.gds374
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.498 15.021 5.538 15.221 ;
 END
 END vccdgt_1p0.gds374
 PIN vccdgt_1p0.gds375
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.458 13.9745 6.498 14.1745 ;
 END
 END vccdgt_1p0.gds375
 PIN vccdgt_1p0.gds376
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.202 13.2695 6.242 13.4695 ;
 END
 END vccdgt_1p0.gds376
 PIN vccdgt_1p0.gds377
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.422 11.9905 7.462 12.1905 ;
 END
 END vccdgt_1p0.gds377
 PIN vccdgt_1p0.gds378
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.67 12.961 6.71 13.161 ;
 END
 END vccdgt_1p0.gds378
 PIN vccdgt_1p0.gds379
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 9.632 15.23 9.688 15.43 ;
 RECT 8.96 15.23 9.016 15.43 ;
 RECT 8.288 15.23 8.344 15.43 ;
 RECT 6.944 15.23 7 15.43 ;
 RECT 7.616 15.23 7.672 15.43 ;
 RECT 9.968 13.197 10.024 13.397 ;
 RECT 9.8 13.197 9.856 13.397 ;
 RECT 10.136 13.197 10.192 13.397 ;
 RECT 9.296 13.197 9.352 13.397 ;
 RECT 9.128 13.197 9.184 13.397 ;
 RECT 9.632 13.214 9.688 13.414 ;
 RECT 9.464 13.197 9.52 13.397 ;
 RECT 8.624 13.197 8.68 13.397 ;
 RECT 8.456 13.197 8.512 13.397 ;
 RECT 8.96 13.214 9.016 13.414 ;
 RECT 8.792 13.197 8.848 13.397 ;
 RECT 7.952 13.197 8.008 13.397 ;
 RECT 7.784 13.197 7.84 13.397 ;
 RECT 8.288 13.214 8.344 13.414 ;
 RECT 8.12 13.197 8.176 13.397 ;
 RECT 7.28 13.197 7.336 13.397 ;
 RECT 7.112 13.197 7.168 13.397 ;
 RECT 6.944 13.214 7 13.414 ;
 RECT 7.616 13.214 7.672 13.414 ;
 RECT 7.448 13.197 7.504 13.397 ;
 RECT 6.272 11.198 6.328 11.398 ;
 RECT 5.348 11.198 5.404 11.398 ;
 RECT 6.104 11.198 6.16 11.398 ;
 RECT 5.852 11.198 5.908 11.398 ;
 RECT 5.684 11.198 5.74 11.398 ;
 RECT 6.44 11.059 6.496 11.259 ;
 RECT 6.44 11.337 6.496 11.537 ;
 RECT 9.968 12.165 10.024 12.365 ;
 RECT 9.8 12.165 9.856 12.365 ;
 RECT 10.136 12.165 10.192 12.365 ;
 RECT 9.296 12.165 9.352 12.365 ;
 RECT 9.128 12.165 9.184 12.365 ;
 RECT 9.464 12.165 9.52 12.365 ;
 RECT 9.632 12.1635 9.688 12.3635 ;
 RECT 8.624 12.165 8.68 12.365 ;
 RECT 8.456 12.165 8.512 12.365 ;
 RECT 8.792 12.165 8.848 12.365 ;
 RECT 8.96 12.1635 9.016 12.3635 ;
 RECT 7.952 12.165 8.008 12.365 ;
 RECT 7.784 12.165 7.84 12.365 ;
 RECT 8.12 12.165 8.176 12.365 ;
 RECT 8.288 12.1635 8.344 12.3635 ;
 RECT 7.28 12.165 7.336 12.365 ;
 RECT 7.112 12.165 7.168 12.365 ;
 RECT 7.448 12.165 7.504 12.365 ;
 RECT 7.616 12.1635 7.672 12.3635 ;
 RECT 6.272 12.542 6.328 12.742 ;
 RECT 5.348 12.542 5.404 12.742 ;
 RECT 6.104 12.542 6.16 12.742 ;
 RECT 5.852 12.542 5.908 12.742 ;
 RECT 6.44 12.403 6.496 12.603 ;
 RECT 5.684 12.542 5.74 12.742 ;
 RECT 6.44 12.681 6.496 12.881 ;
 RECT 5.6 13.886 5.656 14.086 ;
 RECT 5.432 13.886 5.488 14.086 ;
 RECT 5.936 13.886 5.992 14.086 ;
 RECT 5.768 13.886 5.824 14.086 ;
 RECT 6.44 13.886 6.496 14.086 ;
 RECT 6.272 13.886 6.328 14.086 ;
 RECT 6.104 13.886 6.16 14.086 ;
 RECT 5.6 15.23 5.656 15.43 ;
 RECT 5.432 15.23 5.488 15.43 ;
 RECT 5.936 15.23 5.992 15.43 ;
 RECT 5.768 15.23 5.824 15.43 ;
 RECT 6.44 15.23 6.496 15.43 ;
 RECT 6.272 15.23 6.328 15.43 ;
 RECT 6.104 15.23 6.16 15.43 ;
 RECT 6.608 14.8165 6.664 15.0165 ;
 END
 END vccdgt_1p0.gds379
 PIN vccdgt_1p0.gds380
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.422 15.003 13.478 15.203 ;
 END
 END vccdgt_1p0.gds380
 PIN vccdgt_1p0.gds381
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.342 10.662 13.398 10.862 ;
 END
 END vccdgt_1p0.gds381
 PIN vccdgt_1p0.gds382
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.982 11.011 12.042 11.211 ;
 END
 END vccdgt_1p0.gds382
 PIN vccdgt_1p0.gds383
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.814 11.011 11.874 11.211 ;
 END
 END vccdgt_1p0.gds383
 PIN vccdgt_1p0.gds384
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.15 11.011 12.21 11.211 ;
 END
 END vccdgt_1p0.gds384
 PIN vccdgt_1p0.gds385
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.31 11.011 11.37 11.211 ;
 END
 END vccdgt_1p0.gds385
 PIN vccdgt_1p0.gds386
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.142 11.011 11.202 11.211 ;
 END
 END vccdgt_1p0.gds386
 PIN vccdgt_1p0.gds387
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.478 11.011 11.538 11.211 ;
 END
 END vccdgt_1p0.gds387
 PIN vccdgt_1p0.gds388
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.638 11.011 10.698 11.211 ;
 END
 END vccdgt_1p0.gds388
 PIN vccdgt_1p0.gds389
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.47 11.011 10.53 11.211 ;
 END
 END vccdgt_1p0.gds389
 PIN vccdgt_1p0.gds390
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.806 11.011 10.866 11.211 ;
 END
 END vccdgt_1p0.gds390
 PIN vccdgt_1p0.gds391
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.73 12.7505 11.77 12.9505 ;
 END
 END vccdgt_1p0.gds391
 PIN vccdgt_1p0.gds392
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.254 13.309 12.294 13.509 ;
 END
 END vccdgt_1p0.gds392
 PIN vccdgt_1p0.gds393
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.058 12.7505 11.098 12.9505 ;
 END
 END vccdgt_1p0.gds393
 PIN vccdgt_1p0.gds394
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.386 12.7505 10.426 12.9505 ;
 END
 END vccdgt_1p0.gds394
 PIN vccdgt_1p0.gds395
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.186 12.7535 15.226 12.9535 ;
 END
 END vccdgt_1p0.gds395
 PIN vccdgt_1p0.gds396
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.126 11.9905 12.166 12.1905 ;
 END
 END vccdgt_1p0.gds396
 PIN vccdgt_1p0.gds397
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.454 11.9905 11.494 12.1905 ;
 END
 END vccdgt_1p0.gds397
 PIN vccdgt_1p0.gds398
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.782 11.9905 10.822 12.1905 ;
 END
 END vccdgt_1p0.gds398
 PIN vccdgt_1p0.gds399
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.454 15.406 11.494 15.606 ;
 END
 END vccdgt_1p0.gds399
 PIN vccdgt_1p0.gds400
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.782 15.406 10.822 15.606 ;
 END
 END vccdgt_1p0.gds400
 PIN vccdgt_1p0.gds401
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.922 11.224 12.978 11.424 ;
 END
 END vccdgt_1p0.gds401
 PIN vccdgt_1p0.gds402
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.502 10.8945 13.558 11.0945 ;
 END
 END vccdgt_1p0.gds402
 PIN vccdgt_1p0.gds403
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.182 12.7505 14.238 12.9505 ;
 END
 END vccdgt_1p0.gds403
 PIN vccdgt_1p0.gds404
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.766 11.95 14.806 12.15 ;
 END
 END vccdgt_1p0.gds404
 PIN vccdgt_1p0.gds405
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.678 10.478 12.718 10.678 ;
 END
 END vccdgt_1p0.gds405
 PIN vccdgt_1p0.gds406
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.162 13.189 13.238 13.389 ;
 END
 END vccdgt_1p0.gds406
 PIN vccdgt_1p0.gds407
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.922 14.7305 12.978 14.9305 ;
 END
 END vccdgt_1p0.gds407
 PIN vccdgt_1p0.gds408
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.002 13.803 14.078 14.003 ;
 END
 END vccdgt_1p0.gds408
 PIN vccdgt_1p0.gds409
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.126 15.406 12.166 15.606 ;
 END
 END vccdgt_1p0.gds409
 PIN vccdgt_1p0.gds410
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.602 13.638 14.658 13.838 ;
 END
 END vccdgt_1p0.gds410
 PIN vccdgt_1p0.gds411
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.582 13.483 11.622 13.683 ;
 END
 END vccdgt_1p0.gds411
 PIN vccdgt_1p0.gds412
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.934 12.617 11.974 12.817 ;
 END
 END vccdgt_1p0.gds412
 PIN vccdgt_1p0.gds413
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.91 13.483 10.95 13.683 ;
 END
 END vccdgt_1p0.gds413
 PIN vccdgt_1p0.gds414
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.262 12.617 11.302 12.817 ;
 END
 END vccdgt_1p0.gds414
 PIN vccdgt_1p0.gds415
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.238 13.483 10.278 13.683 ;
 END
 END vccdgt_1p0.gds415
 PIN vccdgt_1p0.gds416
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.59 12.617 10.63 12.817 ;
 END
 END vccdgt_1p0.gds416
 PIN vccdgt_1p0.gds417
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.958 14.05 14.998 14.25 ;
 END
 END vccdgt_1p0.gds417
 PIN vccdgt_1p0.gds418
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.402 13.446 12.462 13.646 ;
 END
 END vccdgt_1p0.gds418
 PIN vccdgt_1p0.gds419
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 12.74 15.091 12.796 15.291 ;
 RECT 13.076 15.127 13.132 15.309 ;
 RECT 13.412 15.127 13.468 15.309 ;
 RECT 14.084 15.127 14.14 15.309 ;
 RECT 13.748 15.127 13.804 15.309 ;
 RECT 15.092 15.09 15.148 15.29 ;
 RECT 14.756 15.09 14.812 15.29 ;
 RECT 12.74 15.37 12.796 15.57 ;
 RECT 13.58 15.37 13.636 15.57 ;
 RECT 13.244 15.3035 13.3 15.5035 ;
 RECT 12.908 15.4105 12.964 15.6105 ;
 RECT 13.916 15.2705 13.972 15.4705 ;
 RECT 14.924 15.37 14.98 15.57 ;
 RECT 12.32 15.23 12.376 15.43 ;
 RECT 11.648 15.23 11.704 15.43 ;
 RECT 10.976 15.23 11.032 15.43 ;
 RECT 10.304 15.23 10.36 15.43 ;
 RECT 13.412 14.007 13.468 14.189 ;
 RECT 13.244 13.989 13.3 14.189 ;
 RECT 14.252 14.007 14.308 14.189 ;
 RECT 14.084 14.007 14.14 14.189 ;
 RECT 13.748 14.007 13.804 14.189 ;
 RECT 15.092 14.026 15.148 14.226 ;
 RECT 14.756 14.026 14.812 14.226 ;
 RECT 14.588 14.007 14.644 14.189 ;
 RECT 13.076 13.886 13.132 14.086 ;
 RECT 15.176 13.746 15.232 13.946 ;
 RECT 14.84 13.746 14.896 13.946 ;
 RECT 14.672 13.783 14.728 13.965 ;
 RECT 12.572 14.1515 12.628 14.3515 ;
 RECT 13.496 12.682 13.552 12.882 ;
 RECT 13.076 12.682 13.132 12.882 ;
 RECT 15.176 12.682 15.232 12.882 ;
 RECT 14.84 12.682 14.896 12.882 ;
 RECT 12.656 12.403 12.712 12.603 ;
 RECT 13.412 12.439 13.468 12.621 ;
 RECT 13.244 12.439 13.3 12.621 ;
 RECT 13.076 12.439 13.132 12.621 ;
 RECT 14.336 12.542 14.392 12.742 ;
 RECT 14.084 12.439 14.14 12.621 ;
 RECT 13.916 12.542 13.972 12.742 ;
 RECT 13.748 12.439 13.804 12.621 ;
 RECT 14.84 12.402 14.896 12.602 ;
 RECT 14.672 12.542 14.728 12.742 ;
 RECT 12.656 11.337 12.712 11.537 ;
 RECT 13.076 11.319 13.132 11.501 ;
 RECT 13.412 11.319 13.468 11.501 ;
 RECT 13.244 11.319 13.3 11.501 ;
 RECT 14.336 11.319 14.392 11.501 ;
 RECT 14.084 11.319 14.14 11.501 ;
 RECT 13.916 11.319 13.972 11.501 ;
 RECT 13.748 11.319 13.804 11.501 ;
 RECT 14.84 11.319 14.896 11.501 ;
 RECT 14.672 11.301 14.728 11.501 ;
 RECT 14.924 11.058 14.98 11.258 ;
 RECT 14.588 11.058 14.644 11.258 ;
 RECT 12.908 11.058 12.964 11.258 ;
 RECT 13.916 11.058 13.972 11.258 ;
 RECT 13.58 11.058 13.636 11.258 ;
 RECT 13.244 11.058 13.3 11.258 ;
 RECT 12.656 11.059 12.712 11.259 ;
 RECT 14.252 15.249 14.308 15.449 ;
 RECT 14.252 10.988 14.308 11.188 ;
 RECT 11.984 13.197 12.04 13.397 ;
 RECT 11.816 13.197 11.872 13.397 ;
 RECT 12.32 13.214 12.376 13.414 ;
 RECT 12.152 13.197 12.208 13.397 ;
 RECT 11.312 13.197 11.368 13.397 ;
 RECT 11.144 13.197 11.2 13.397 ;
 RECT 11.648 13.214 11.704 13.414 ;
 RECT 11.48 13.197 11.536 13.397 ;
 RECT 10.64 13.197 10.696 13.397 ;
 RECT 10.472 13.197 10.528 13.397 ;
 RECT 10.976 13.214 11.032 13.414 ;
 RECT 10.808 13.197 10.864 13.397 ;
 RECT 10.304 13.214 10.36 13.414 ;
 RECT 12.908 13.634 12.964 13.834 ;
 RECT 13.496 13.676 13.552 13.876 ;
 RECT 13.916 13.7925 13.972 13.9925 ;
 RECT 14.336 13.676 14.392 13.876 ;
 RECT 14.504 15.2025 14.56 15.4025 ;
 RECT 11.984 12.165 12.04 12.365 ;
 RECT 11.816 12.165 11.872 12.365 ;
 RECT 12.152 12.165 12.208 12.365 ;
 RECT 12.32 12.1635 12.376 12.3635 ;
 RECT 11.312 12.165 11.368 12.365 ;
 RECT 11.144 12.165 11.2 12.365 ;
 RECT 11.48 12.165 11.536 12.365 ;
 RECT 11.648 12.1635 11.704 12.3635 ;
 RECT 10.64 12.165 10.696 12.365 ;
 RECT 10.472 12.165 10.528 12.365 ;
 RECT 10.808 12.165 10.864 12.365 ;
 RECT 10.976 12.1635 11.032 12.3635 ;
 RECT 10.304 12.1635 10.36 12.3635 ;
 END
 END vccdgt_1p0.gds419
 PIN vccdgt_1p0.gds420
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.626 12.7505 19.666 12.9505 ;
 END
 END vccdgt_1p0.gds420
 PIN vccdgt_1p0.gds421
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.71 11.011 19.77 11.211 ;
 END
 END vccdgt_1p0.gds421
 PIN vccdgt_1p0.gds422
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.038 11.011 19.098 11.211 ;
 END
 END vccdgt_1p0.gds422
 PIN vccdgt_1p0.gds423
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.366 11.011 18.426 11.211 ;
 END
 END vccdgt_1p0.gds423
 PIN vccdgt_1p0.gds424
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 10.502 16.57 10.702 ;
 END
 END vccdgt_1p0.gds424
 PIN vccdgt_1p0.gds425
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.838 12.5175 16.894 12.7175 ;
 END
 END vccdgt_1p0.gds425
 PIN vccdgt_1p0.gds426
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.878 11.011 19.938 11.211 ;
 END
 END vccdgt_1p0.gds426
 PIN vccdgt_1p0.gds427
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.046 11.011 20.106 11.211 ;
 END
 END vccdgt_1p0.gds427
 PIN vccdgt_1p0.gds428
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.206 11.011 19.266 11.211 ;
 END
 END vccdgt_1p0.gds428
 PIN vccdgt_1p0.gds429
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.374 11.011 19.434 11.211 ;
 END
 END vccdgt_1p0.gds429
 PIN vccdgt_1p0.gds430
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.534 11.011 18.594 11.211 ;
 END
 END vccdgt_1p0.gds430
 PIN vccdgt_1p0.gds431
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.702 11.011 18.762 11.211 ;
 END
 END vccdgt_1p0.gds431
 PIN vccdgt_1p0.gds432
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.866 14.062 15.926 14.262 ;
 END
 END vccdgt_1p0.gds432
 PIN vccdgt_1p0.gds433
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.018 13.1425 17.074 13.3425 ;
 END
 END vccdgt_1p0.gds433
 PIN vccdgt_1p0.gds434
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.954 12.7505 18.994 12.9505 ;
 END
 END vccdgt_1p0.gds434
 PIN vccdgt_1p0.gds435
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.282 12.7505 18.322 12.9505 ;
 END
 END vccdgt_1p0.gds435
 PIN vccdgt_1p0.gds436
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.022 15.406 20.062 15.606 ;
 END
 END vccdgt_1p0.gds436
 PIN vccdgt_1p0.gds437
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.35 15.406 19.39 15.606 ;
 END
 END vccdgt_1p0.gds437
 PIN vccdgt_1p0.gds438
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.022 11.9905 20.062 12.1905 ;
 END
 END vccdgt_1p0.gds438
 PIN vccdgt_1p0.gds439
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.15 13.483 20.19 13.683 ;
 END
 END vccdgt_1p0.gds439
 PIN vccdgt_1p0.gds440
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.478 13.483 19.518 13.683 ;
 END
 END vccdgt_1p0.gds440
 PIN vccdgt_1p0.gds441
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.83 12.617 19.87 12.817 ;
 END
 END vccdgt_1p0.gds441
 PIN vccdgt_1p0.gds442
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.03 14.161 16.076 14.361 ;
 END
 END vccdgt_1p0.gds442
 PIN vccdgt_1p0.gds443
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 13.374 17.734 13.574 ;
 END
 END vccdgt_1p0.gds443
 PIN vccdgt_1p0.gds444
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.314 13.2495 15.354 13.4495 ;
 END
 END vccdgt_1p0.gds444
 PIN vccdgt_1p0.gds445
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.334 13.268 16.39 13.468 ;
 END
 END vccdgt_1p0.gds445
 PIN vccdgt_1p0.gds446
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.338 13.2505 17.414 13.4505 ;
 END
 END vccdgt_1p0.gds446
 PIN vccdgt_1p0.gds447
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.522 12.3155 15.582 12.5155 ;
 END
 END vccdgt_1p0.gds447
 PIN vccdgt_1p0.gds448
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.598 11.025 17.654 11.225 ;
 END
 END vccdgt_1p0.gds448
 PIN vccdgt_1p0.gds449
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.674 12.968 16.734 13.168 ;
 END
 END vccdgt_1p0.gds449
 PIN vccdgt_1p0.gds450
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.858 11.6505 17.898 11.8505 ;
 END
 END vccdgt_1p0.gds450
 PIN vccdgt_1p0.gds451
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.158 12.617 19.198 12.817 ;
 END
 END vccdgt_1p0.gds451
 PIN vccdgt_1p0.gds452
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.486 12.617 18.526 12.817 ;
 END
 END vccdgt_1p0.gds452
 PIN vccdgt_1p0.gds453
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.806 13.483 18.846 13.683 ;
 END
 END vccdgt_1p0.gds453
 PIN vccdgt_1p0.gds454
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.35 11.9905 19.39 12.1905 ;
 END
 END vccdgt_1p0.gds454
 PIN vccdgt_1p0.gds455
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.678 11.9905 18.718 12.1905 ;
 END
 END vccdgt_1p0.gds455
 PIN vccdgt_1p0.gds456
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.114 13.2825 18.174 13.4825 ;
 END
 END vccdgt_1p0.gds456
 PIN vccdgt_1p0.gds457
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.178 13.0715 17.234 13.2715 ;
 END
 END vccdgt_1p0.gds457
 PIN vccdgt_1p0.gds458
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.678 15.406 18.718 15.606 ;
 END
 END vccdgt_1p0.gds458
 PIN vccdgt_1p0.gds459
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 15.428 15.09 15.484 15.29 ;
 RECT 16.688 15.109 16.744 15.309 ;
 RECT 16.268 15.127 16.324 15.309 ;
 RECT 17.78 15.091 17.836 15.291 ;
 RECT 20.216 15.23 20.272 15.43 ;
 RECT 15.26 15.37 15.316 15.57 ;
 RECT 15.932 15.37 15.988 15.57 ;
 RECT 15.596 15.37 15.652 15.57 ;
 RECT 16.268 15.37 16.324 15.57 ;
 RECT 17.528 15.23 17.584 15.43 ;
 RECT 17.192 15.351 17.248 15.533 ;
 RECT 17.78 15.369 17.836 15.569 ;
 RECT 19.544 15.23 19.6 15.43 ;
 RECT 18.2 15.23 18.256 15.43 ;
 RECT 18.872 15.23 18.928 15.43 ;
 RECT 15.512 13.746 15.568 13.946 ;
 RECT 15.848 13.785 15.904 13.951 ;
 RECT 16.1 12.679 16.156 12.843 ;
 RECT 15.512 12.682 15.568 12.882 ;
 RECT 15.848 12.672 15.904 12.843 ;
 RECT 17.528 12.681 17.584 12.881 ;
 RECT 15.932 12.439 15.988 12.621 ;
 RECT 15.764 12.439 15.82 12.621 ;
 RECT 15.596 12.439 15.652 12.621 ;
 RECT 15.428 12.439 15.484 12.621 ;
 RECT 16.604 12.403 16.66 12.603 ;
 RECT 16.184 12.441 16.24 12.621 ;
 RECT 17.528 12.403 17.584 12.603 ;
 RECT 16.94 12.402 16.996 12.602 ;
 RECT 17.78 12.403 17.836 12.603 ;
 RECT 15.764 11.301 15.82 11.501 ;
 RECT 15.596 11.301 15.652 11.501 ;
 RECT 15.428 11.301 15.484 11.501 ;
 RECT 16.688 11.338 16.744 11.538 ;
 RECT 16.52 11.301 16.576 11.501 ;
 RECT 16.352 11.301 16.408 11.501 ;
 RECT 17.528 11.301 17.584 11.501 ;
 RECT 17.864 11.337 17.92 11.537 ;
 RECT 16.604 11.058 16.66 11.258 ;
 RECT 16.94 11.058 16.996 11.258 ;
 RECT 17.108 12.3615 17.164 12.5615 ;
 RECT 17.276 12.3615 17.332 12.5615 ;
 RECT 16.268 10.988 16.324 11.188 ;
 RECT 15.932 11.1275 15.988 11.3275 ;
 RECT 16.184 11.2685 16.24 11.4685 ;
 RECT 18.032 14.5165 18.088 14.7165 ;
 RECT 17.024 12.752 17.08 12.952 ;
 RECT 16.52 12.752 16.576 12.952 ;
 RECT 19.88 13.197 19.936 13.397 ;
 RECT 19.712 13.197 19.768 13.397 ;
 RECT 20.216 13.214 20.272 13.414 ;
 RECT 20.048 13.197 20.104 13.397 ;
 RECT 19.208 13.197 19.264 13.397 ;
 RECT 19.04 13.197 19.096 13.397 ;
 RECT 19.544 13.214 19.6 13.414 ;
 RECT 19.376 13.197 19.432 13.397 ;
 RECT 18.536 13.197 18.592 13.397 ;
 RECT 18.368 13.197 18.424 13.397 ;
 RECT 18.2 13.214 18.256 13.414 ;
 RECT 18.872 13.214 18.928 13.414 ;
 RECT 18.704 13.197 18.76 13.397 ;
 RECT 19.88 12.165 19.936 12.365 ;
 RECT 19.712 12.165 19.768 12.365 ;
 RECT 20.048 12.165 20.104 12.365 ;
 RECT 20.216 12.1635 20.272 12.3635 ;
 RECT 19.208 12.165 19.264 12.365 ;
 RECT 19.04 12.165 19.096 12.365 ;
 RECT 19.376 12.165 19.432 12.365 ;
 RECT 19.544 12.1635 19.6 12.3635 ;
 RECT 18.536 12.165 18.592 12.365 ;
 RECT 18.368 12.165 18.424 12.365 ;
 RECT 18.704 12.165 18.76 12.365 ;
 RECT 18.872 12.1635 18.928 12.3635 ;
 RECT 15.848 15.02 15.904 15.22 ;
 RECT 17.276 15.02 17.332 15.22 ;
 RECT 17.108 15.02 17.164 15.22 ;
 RECT 16.016 15.09 16.072 15.29 ;
 RECT 16.52 15.127 16.576 15.309 ;
 RECT 17.444 15.239 17.5 15.439 ;
 RECT 16.94 15.351 16.996 15.533 ;
 RECT 17.696 11.267 17.752 11.467 ;
 RECT 16.94 11.408 16.996 11.608 ;
 RECT 17.108 11.408 17.164 11.608 ;
 RECT 17.276 11.291 17.332 11.491 ;
 RECT 16.604 13.676 16.66 13.876 ;
 RECT 17.528 13.7265 17.584 13.9265 ;
 RECT 17.108 13.676 17.164 13.876 ;
 RECT 16.1 13.8845 16.156 14.0845 ;
 RECT 15.428 14.026 15.484 14.226 ;
 RECT 15.932 14.007 15.988 14.189 ;
 RECT 15.764 14.007 15.82 14.189 ;
 RECT 16.688 14.007 16.744 14.189 ;
 RECT 16.52 14.007 16.576 14.189 ;
 RECT 16.352 14.007 16.408 14.189 ;
 RECT 17.36 14.007 17.416 14.189 ;
 RECT 17.192 14.007 17.248 14.189 ;
 RECT 18.116 14.064 18.172 14.264 ;
 END
 END vccdgt_1p0.gds459
 PIN vccdgt_1p0.gds460
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.078 12.7505 24.118 12.9505 ;
 END
 END vccdgt_1p0.gds460
 PIN vccdgt_1p0.gds461
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.986 12.7505 23.026 12.9505 ;
 END
 END vccdgt_1p0.gds461
 PIN vccdgt_1p0.gds462
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.75 12.7505 24.79 12.9505 ;
 END
 END vccdgt_1p0.gds462
 PIN vccdgt_1p0.gds463
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.51 13.309 23.55 13.509 ;
 END
 END vccdgt_1p0.gds463
 PIN vccdgt_1p0.gds464
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.314 12.7505 22.354 12.9505 ;
 END
 END vccdgt_1p0.gds464
 PIN vccdgt_1p0.gds465
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.642 12.7505 21.682 12.9505 ;
 END
 END vccdgt_1p0.gds465
 PIN vccdgt_1p0.gds466
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.97 12.7505 21.01 12.9505 ;
 END
 END vccdgt_1p0.gds466
 PIN vccdgt_1p0.gds467
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.298 12.7505 20.338 12.9505 ;
 END
 END vccdgt_1p0.gds467
 PIN vccdgt_1p0.gds468
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.834 11.011 24.894 11.211 ;
 END
 END vccdgt_1p0.gds468
 PIN vccdgt_1p0.gds469
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.162 11.011 24.222 11.211 ;
 END
 END vccdgt_1p0.gds469
 PIN vccdgt_1p0.gds470
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.07 11.011 23.13 11.211 ;
 END
 END vccdgt_1p0.gds470
 PIN vccdgt_1p0.gds471
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.398 11.011 22.458 11.211 ;
 END
 END vccdgt_1p0.gds471
 PIN vccdgt_1p0.gds472
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.726 11.011 21.786 11.211 ;
 END
 END vccdgt_1p0.gds472
 PIN vccdgt_1p0.gds473
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.054 11.011 21.114 11.211 ;
 END
 END vccdgt_1p0.gds473
 PIN vccdgt_1p0.gds474
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.382 11.011 20.442 11.211 ;
 END
 END vccdgt_1p0.gds474
 PIN vccdgt_1p0.gds475
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.002 11.011 25.062 11.211 ;
 END
 END vccdgt_1p0.gds475
 PIN vccdgt_1p0.gds476
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.17 11.011 25.23 11.211 ;
 END
 END vccdgt_1p0.gds476
 PIN vccdgt_1p0.gds477
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.33 11.011 24.39 11.211 ;
 END
 END vccdgt_1p0.gds477
 PIN vccdgt_1p0.gds478
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.498 11.011 24.558 11.211 ;
 END
 END vccdgt_1p0.gds478
 PIN vccdgt_1p0.gds479
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.238 11.011 23.298 11.211 ;
 END
 END vccdgt_1p0.gds479
 PIN vccdgt_1p0.gds480
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.406 11.011 23.466 11.211 ;
 END
 END vccdgt_1p0.gds480
 PIN vccdgt_1p0.gds481
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.566 11.011 22.626 11.211 ;
 END
 END vccdgt_1p0.gds481
 PIN vccdgt_1p0.gds482
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.734 11.011 22.794 11.211 ;
 END
 END vccdgt_1p0.gds482
 PIN vccdgt_1p0.gds483
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.894 11.011 21.954 11.211 ;
 END
 END vccdgt_1p0.gds483
 PIN vccdgt_1p0.gds484
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.062 11.011 22.122 11.211 ;
 END
 END vccdgt_1p0.gds484
 PIN vccdgt_1p0.gds485
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.222 11.011 21.282 11.211 ;
 END
 END vccdgt_1p0.gds485
 PIN vccdgt_1p0.gds486
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.39 11.011 21.45 11.211 ;
 END
 END vccdgt_1p0.gds486
 PIN vccdgt_1p0.gds487
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.55 11.011 20.61 11.211 ;
 END
 END vccdgt_1p0.gds487
 PIN vccdgt_1p0.gds488
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.718 11.011 20.778 11.211 ;
 END
 END vccdgt_1p0.gds488
 PIN vccdgt_1p0.gds489
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.146 15.406 25.186 15.606 ;
 END
 END vccdgt_1p0.gds489
 PIN vccdgt_1p0.gds490
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.71 15.406 22.75 15.606 ;
 END
 END vccdgt_1p0.gds490
 PIN vccdgt_1p0.gds491
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.038 15.406 22.078 15.606 ;
 END
 END vccdgt_1p0.gds491
 PIN vccdgt_1p0.gds492
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.366 15.406 21.406 15.606 ;
 END
 END vccdgt_1p0.gds492
 PIN vccdgt_1p0.gds493
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.694 15.406 20.734 15.606 ;
 END
 END vccdgt_1p0.gds493
 PIN vccdgt_1p0.gds494
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.146 11.9905 25.186 12.1905 ;
 END
 END vccdgt_1p0.gds494
 PIN vccdgt_1p0.gds495
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.474 11.9905 24.514 12.1905 ;
 END
 END vccdgt_1p0.gds495
 PIN vccdgt_1p0.gds496
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.382 11.9905 23.422 12.1905 ;
 END
 END vccdgt_1p0.gds496
 PIN vccdgt_1p0.gds497
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.71 11.9905 22.75 12.1905 ;
 END
 END vccdgt_1p0.gds497
 PIN vccdgt_1p0.gds498
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.038 11.9905 22.078 12.1905 ;
 END
 END vccdgt_1p0.gds498
 PIN vccdgt_1p0.gds499
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.366 11.9905 21.406 12.1905 ;
 END
 END vccdgt_1p0.gds499
 PIN vccdgt_1p0.gds500
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.694 11.9905 20.734 12.1905 ;
 END
 END vccdgt_1p0.gds500
 PIN vccdgt_1p0.gds501
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.602 13.483 24.642 13.683 ;
 END
 END vccdgt_1p0.gds501
 PIN vccdgt_1p0.gds502
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.954 12.617 24.994 12.817 ;
 END
 END vccdgt_1p0.gds502
 PIN vccdgt_1p0.gds503
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.93 13.4245 23.97 13.6245 ;
 END
 END vccdgt_1p0.gds503
 PIN vccdgt_1p0.gds504
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.282 12.617 24.322 12.817 ;
 END
 END vccdgt_1p0.gds504
 PIN vccdgt_1p0.gds505
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.838 13.483 22.878 13.683 ;
 END
 END vccdgt_1p0.gds505
 PIN vccdgt_1p0.gds506
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.19 12.617 23.23 12.817 ;
 END
 END vccdgt_1p0.gds506
 PIN vccdgt_1p0.gds507
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.166 13.483 22.206 13.683 ;
 END
 END vccdgt_1p0.gds507
 PIN vccdgt_1p0.gds508
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.518 12.617 22.558 12.817 ;
 END
 END vccdgt_1p0.gds508
 PIN vccdgt_1p0.gds509
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.494 13.483 21.534 13.683 ;
 END
 END vccdgt_1p0.gds509
 PIN vccdgt_1p0.gds510
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.846 12.617 21.886 12.817 ;
 END
 END vccdgt_1p0.gds510
 PIN vccdgt_1p0.gds511
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.822 13.483 20.862 13.683 ;
 END
 END vccdgt_1p0.gds511
 PIN vccdgt_1p0.gds512
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.174 12.617 21.214 12.817 ;
 END
 END vccdgt_1p0.gds512
 PIN vccdgt_1p0.gds513
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.502 12.617 20.542 12.817 ;
 END
 END vccdgt_1p0.gds513
 PIN vccdgt_1p0.gds514
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.474 15.406 24.514 15.606 ;
 END
 END vccdgt_1p0.gds514
 PIN vccdgt_1p0.gds515
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.382 15.406 23.422 15.606 ;
 END
 END vccdgt_1p0.gds515
 PIN vccdgt_1p0.gds516
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.658 13.0135 23.698 13.2135 ;
 END
 END vccdgt_1p0.gds516
 PIN vccdgt_1p0.gds517
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 23.996 15.23 24.052 15.43 ;
 RECT 24.668 15.23 24.724 15.43 ;
 RECT 23.576 15.23 23.632 15.43 ;
 RECT 22.904 15.23 22.96 15.43 ;
 RECT 22.232 15.23 22.288 15.43 ;
 RECT 21.56 15.23 21.616 15.43 ;
 RECT 20.888 15.23 20.944 15.43 ;
 RECT 25.004 13.197 25.06 13.397 ;
 RECT 24.836 13.197 24.892 13.397 ;
 RECT 25.172 13.197 25.228 13.397 ;
 RECT 24.332 13.197 24.388 13.397 ;
 RECT 24.164 13.197 24.22 13.397 ;
 RECT 23.996 13.214 24.052 13.414 ;
 RECT 24.668 13.214 24.724 13.414 ;
 RECT 24.5 13.197 24.556 13.397 ;
 RECT 23.24 13.197 23.296 13.397 ;
 RECT 23.072 13.197 23.128 13.397 ;
 RECT 23.576 13.214 23.632 13.414 ;
 RECT 23.408 13.197 23.464 13.397 ;
 RECT 22.568 13.197 22.624 13.397 ;
 RECT 22.4 13.197 22.456 13.397 ;
 RECT 22.904 13.214 22.96 13.414 ;
 RECT 22.736 13.197 22.792 13.397 ;
 RECT 21.896 13.197 21.952 13.397 ;
 RECT 21.728 13.197 21.784 13.397 ;
 RECT 22.232 13.214 22.288 13.414 ;
 RECT 22.064 13.197 22.12 13.397 ;
 RECT 21.224 13.197 21.28 13.397 ;
 RECT 21.056 13.197 21.112 13.397 ;
 RECT 21.56 13.214 21.616 13.414 ;
 RECT 21.392 13.197 21.448 13.397 ;
 RECT 20.552 13.197 20.608 13.397 ;
 RECT 20.888 13.214 20.944 13.414 ;
 RECT 20.72 13.197 20.776 13.397 ;
 RECT 20.384 13.197 20.44 13.397 ;
 RECT 25.004 12.165 25.06 12.365 ;
 RECT 24.836 12.165 24.892 12.365 ;
 RECT 25.172 12.165 25.228 12.365 ;
 RECT 24.332 12.165 24.388 12.365 ;
 RECT 24.164 12.165 24.22 12.365 ;
 RECT 24.5 12.165 24.556 12.365 ;
 RECT 24.668 12.1635 24.724 12.3635 ;
 RECT 23.24 12.165 23.296 12.365 ;
 RECT 23.072 12.165 23.128 12.365 ;
 RECT 23.408 12.165 23.464 12.365 ;
 RECT 23.576 12.1635 23.632 12.3635 ;
 RECT 22.568 12.165 22.624 12.365 ;
 RECT 22.4 12.165 22.456 12.365 ;
 RECT 22.736 12.165 22.792 12.365 ;
 RECT 22.904 12.1635 22.96 12.3635 ;
 RECT 21.896 12.165 21.952 12.365 ;
 RECT 21.728 12.165 21.784 12.365 ;
 RECT 22.064 12.165 22.12 12.365 ;
 RECT 22.232 12.1635 22.288 12.3635 ;
 RECT 21.224 12.165 21.28 12.365 ;
 RECT 21.056 12.165 21.112 12.365 ;
 RECT 21.392 12.165 21.448 12.365 ;
 RECT 21.56 12.1635 21.616 12.3635 ;
 RECT 20.552 12.165 20.608 12.365 ;
 RECT 20.72 12.165 20.776 12.365 ;
 RECT 20.888 12.1635 20.944 12.3635 ;
 RECT 20.384 12.165 20.44 12.365 ;
 RECT 23.828 13.659 23.884 13.859 ;
 RECT 23.912 13.095 23.968 13.295 ;
 RECT 23.66 13.2495 23.716 13.4495 ;
 END
 END vccdgt_1p0.gds517
 PIN vccdgt_1p0.gds518
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.782 12.7505 28.822 12.9505 ;
 END
 END vccdgt_1p0.gds518
 PIN vccdgt_1p0.gds519
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.306 13.309 29.346 13.509 ;
 END
 END vccdgt_1p0.gds519
 PIN vccdgt_1p0.gds520
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.11 12.7505 28.15 12.9505 ;
 END
 END vccdgt_1p0.gds520
 PIN vccdgt_1p0.gds521
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.438 12.7505 27.478 12.9505 ;
 END
 END vccdgt_1p0.gds521
 PIN vccdgt_1p0.gds522
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.766 12.7505 26.806 12.9505 ;
 END
 END vccdgt_1p0.gds522
 PIN vccdgt_1p0.gds523
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.094 12.7505 26.134 12.9505 ;
 END
 END vccdgt_1p0.gds523
 PIN vccdgt_1p0.gds524
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.422 12.7505 25.462 12.9505 ;
 END
 END vccdgt_1p0.gds524
 PIN vccdgt_1p0.gds525
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.866 11.011 28.926 11.211 ;
 END
 END vccdgt_1p0.gds525
 PIN vccdgt_1p0.gds526
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.194 11.011 28.254 11.211 ;
 END
 END vccdgt_1p0.gds526
 PIN vccdgt_1p0.gds527
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.522 11.011 27.582 11.211 ;
 END
 END vccdgt_1p0.gds527
 PIN vccdgt_1p0.gds528
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.85 11.011 26.91 11.211 ;
 END
 END vccdgt_1p0.gds528
 PIN vccdgt_1p0.gds529
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.178 11.011 26.238 11.211 ;
 END
 END vccdgt_1p0.gds529
 PIN vccdgt_1p0.gds530
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.506 11.011 25.566 11.211 ;
 END
 END vccdgt_1p0.gds530
 PIN vccdgt_1p0.gds531
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.034 11.011 29.094 11.211 ;
 END
 END vccdgt_1p0.gds531
 PIN vccdgt_1p0.gds532
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.202 11.011 29.262 11.211 ;
 END
 END vccdgt_1p0.gds532
 PIN vccdgt_1p0.gds533
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.362 11.011 28.422 11.211 ;
 END
 END vccdgt_1p0.gds533
 PIN vccdgt_1p0.gds534
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.53 11.011 28.59 11.211 ;
 END
 END vccdgt_1p0.gds534
 PIN vccdgt_1p0.gds535
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.69 11.011 27.75 11.211 ;
 END
 END vccdgt_1p0.gds535
 PIN vccdgt_1p0.gds536
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.858 11.011 27.918 11.211 ;
 END
 END vccdgt_1p0.gds536
 PIN vccdgt_1p0.gds537
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.018 11.011 27.078 11.211 ;
 END
 END vccdgt_1p0.gds537
 PIN vccdgt_1p0.gds538
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.186 11.011 27.246 11.211 ;
 END
 END vccdgt_1p0.gds538
 PIN vccdgt_1p0.gds539
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.346 11.011 26.406 11.211 ;
 END
 END vccdgt_1p0.gds539
 PIN vccdgt_1p0.gds540
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.514 11.011 26.574 11.211 ;
 END
 END vccdgt_1p0.gds540
 PIN vccdgt_1p0.gds541
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.674 11.011 25.734 11.211 ;
 END
 END vccdgt_1p0.gds541
 PIN vccdgt_1p0.gds542
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.842 11.011 25.902 11.211 ;
 END
 END vccdgt_1p0.gds542
 PIN vccdgt_1p0.gds543
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.506 15.406 28.546 15.606 ;
 END
 END vccdgt_1p0.gds543
 PIN vccdgt_1p0.gds544
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.834 15.406 27.874 15.606 ;
 END
 END vccdgt_1p0.gds544
 PIN vccdgt_1p0.gds545
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.162 15.406 27.202 15.606 ;
 END
 END vccdgt_1p0.gds545
 PIN vccdgt_1p0.gds546
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.49 15.406 26.53 15.606 ;
 END
 END vccdgt_1p0.gds546
 PIN vccdgt_1p0.gds547
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.818 15.406 25.858 15.606 ;
 END
 END vccdgt_1p0.gds547
 PIN vccdgt_1p0.gds548
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.178 11.9905 29.218 12.1905 ;
 END
 END vccdgt_1p0.gds548
 PIN vccdgt_1p0.gds549
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.506 11.9905 28.546 12.1905 ;
 END
 END vccdgt_1p0.gds549
 PIN vccdgt_1p0.gds550
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.834 11.9905 27.874 12.1905 ;
 END
 END vccdgt_1p0.gds550
 PIN vccdgt_1p0.gds551
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.162 11.9905 27.202 12.1905 ;
 END
 END vccdgt_1p0.gds551
 PIN vccdgt_1p0.gds552
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.49 11.9905 26.53 12.1905 ;
 END
 END vccdgt_1p0.gds552
 PIN vccdgt_1p0.gds553
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.818 11.9905 25.858 12.1905 ;
 END
 END vccdgt_1p0.gds553
 PIN vccdgt_1p0.gds554
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.634 13.483 28.674 13.683 ;
 END
 END vccdgt_1p0.gds554
 PIN vccdgt_1p0.gds555
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.986 12.617 29.026 12.817 ;
 END
 END vccdgt_1p0.gds555
 PIN vccdgt_1p0.gds556
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.962 13.483 28.002 13.683 ;
 END
 END vccdgt_1p0.gds556
 PIN vccdgt_1p0.gds557
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.314 12.617 28.354 12.817 ;
 END
 END vccdgt_1p0.gds557
 PIN vccdgt_1p0.gds558
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.29 13.483 27.33 13.683 ;
 END
 END vccdgt_1p0.gds558
 PIN vccdgt_1p0.gds559
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.642 12.617 27.682 12.817 ;
 END
 END vccdgt_1p0.gds559
 PIN vccdgt_1p0.gds560
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.618 13.483 26.658 13.683 ;
 END
 END vccdgt_1p0.gds560
 PIN vccdgt_1p0.gds561
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.97 12.617 27.01 12.817 ;
 END
 END vccdgt_1p0.gds561
 PIN vccdgt_1p0.gds562
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.946 13.483 25.986 13.683 ;
 END
 END vccdgt_1p0.gds562
 PIN vccdgt_1p0.gds563
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.298 12.617 26.338 12.817 ;
 END
 END vccdgt_1p0.gds563
 PIN vccdgt_1p0.gds564
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.274 13.483 25.314 13.683 ;
 END
 END vccdgt_1p0.gds564
 PIN vccdgt_1p0.gds565
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.626 12.617 25.666 12.817 ;
 END
 END vccdgt_1p0.gds565
 PIN vccdgt_1p0.gds566
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.974 14.7305 30.03 14.9305 ;
 END
 END vccdgt_1p0.gds566
 PIN vccdgt_1p0.gds567
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.178 15.406 29.218 15.606 ;
 END
 END vccdgt_1p0.gds567
 PIN vccdgt_1p0.gds568
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.214 13.189 30.29 13.389 ;
 END
 END vccdgt_1p0.gds568
 PIN vccdgt_1p0.gds569
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.974 11.224 30.03 11.424 ;
 END
 END vccdgt_1p0.gds569
 PIN vccdgt_1p0.gds570
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.73 10.478 29.77 10.678 ;
 END
 END vccdgt_1p0.gds570
 PIN vccdgt_1p0.gds571
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.454 13.446 29.514 13.646 ;
 END
 END vccdgt_1p0.gds571
 PIN vccdgt_1p0.gds572
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 29.792 15.091 29.848 15.291 ;
 RECT 30.128 15.127 30.184 15.309 ;
 RECT 29.792 15.37 29.848 15.57 ;
 RECT 29.96 15.4105 30.016 15.6105 ;
 RECT 29.372 15.23 29.428 15.43 ;
 RECT 28.7 15.23 28.756 15.43 ;
 RECT 28.028 15.23 28.084 15.43 ;
 RECT 27.356 15.23 27.412 15.43 ;
 RECT 26.684 15.23 26.74 15.43 ;
 RECT 26.012 15.23 26.068 15.43 ;
 RECT 25.34 15.23 25.396 15.43 ;
 RECT 30.128 12.682 30.184 12.882 ;
 RECT 29.708 12.403 29.764 12.603 ;
 RECT 30.128 12.439 30.184 12.621 ;
 RECT 29.708 11.337 29.764 11.537 ;
 RECT 30.128 11.319 30.184 11.501 ;
 RECT 29.96 11.058 30.016 11.258 ;
 RECT 29.708 11.059 29.764 11.259 ;
 RECT 29.96 13.634 30.016 13.834 ;
 RECT 30.128 13.886 30.184 14.086 ;
 RECT 29.624 14.1515 29.68 14.3515 ;
 RECT 29.036 13.197 29.092 13.397 ;
 RECT 28.868 13.197 28.924 13.397 ;
 RECT 29.372 13.214 29.428 13.414 ;
 RECT 29.204 13.197 29.26 13.397 ;
 RECT 28.364 13.197 28.42 13.397 ;
 RECT 28.196 13.197 28.252 13.397 ;
 RECT 28.7 13.214 28.756 13.414 ;
 RECT 28.532 13.197 28.588 13.397 ;
 RECT 27.692 13.197 27.748 13.397 ;
 RECT 27.524 13.197 27.58 13.397 ;
 RECT 28.028 13.214 28.084 13.414 ;
 RECT 27.86 13.197 27.916 13.397 ;
 RECT 27.02 13.197 27.076 13.397 ;
 RECT 26.852 13.197 26.908 13.397 ;
 RECT 27.356 13.214 27.412 13.414 ;
 RECT 27.188 13.197 27.244 13.397 ;
 RECT 26.348 13.197 26.404 13.397 ;
 RECT 26.18 13.197 26.236 13.397 ;
 RECT 26.684 13.214 26.74 13.414 ;
 RECT 26.516 13.197 26.572 13.397 ;
 RECT 25.676 13.197 25.732 13.397 ;
 RECT 25.508 13.197 25.564 13.397 ;
 RECT 26.012 13.214 26.068 13.414 ;
 RECT 25.844 13.197 25.9 13.397 ;
 RECT 25.34 13.214 25.396 13.414 ;
 RECT 29.036 12.165 29.092 12.365 ;
 RECT 28.868 12.165 28.924 12.365 ;
 RECT 29.204 12.165 29.26 12.365 ;
 RECT 29.372 12.1635 29.428 12.3635 ;
 RECT 28.364 12.165 28.42 12.365 ;
 RECT 28.196 12.165 28.252 12.365 ;
 RECT 28.532 12.165 28.588 12.365 ;
 RECT 28.7 12.1635 28.756 12.3635 ;
 RECT 27.692 12.165 27.748 12.365 ;
 RECT 27.524 12.165 27.58 12.365 ;
 RECT 27.86 12.165 27.916 12.365 ;
 RECT 28.028 12.1635 28.084 12.3635 ;
 RECT 27.02 12.165 27.076 12.365 ;
 RECT 26.852 12.165 26.908 12.365 ;
 RECT 27.188 12.165 27.244 12.365 ;
 RECT 27.356 12.1635 27.412 12.3635 ;
 RECT 26.348 12.165 26.404 12.365 ;
 RECT 26.18 12.165 26.236 12.365 ;
 RECT 26.516 12.165 26.572 12.365 ;
 RECT 26.684 12.1635 26.74 12.3635 ;
 RECT 25.676 12.165 25.732 12.365 ;
 RECT 25.508 12.165 25.564 12.365 ;
 RECT 25.844 12.165 25.9 12.365 ;
 RECT 26.012 12.1635 26.068 12.3635 ;
 RECT 25.34 12.1635 25.396 12.3635 ;
 END
 END vccdgt_1p0.gds572
 PIN vccdgt_1p0.gds573
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.07 13.1425 34.126 13.3425 ;
 END
 END vccdgt_1p0.gds573
 PIN vccdgt_1p0.gds574
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.474 15.003 30.53 15.203 ;
 END
 END vccdgt_1p0.gds574
 PIN vccdgt_1p0.gds575
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 10.502 33.622 10.702 ;
 END
 END vccdgt_1p0.gds575
 PIN vccdgt_1p0.gds576
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.89 12.5175 33.946 12.7175 ;
 END
 END vccdgt_1p0.gds576
 PIN vccdgt_1p0.gds577
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.918 14.062 32.978 14.262 ;
 END
 END vccdgt_1p0.gds577
 PIN vccdgt_1p0.gds578
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.394 10.662 30.45 10.862 ;
 END
 END vccdgt_1p0.gds578
 PIN vccdgt_1p0.gds579
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.39 13.2505 34.466 13.4505 ;
 END
 END vccdgt_1p0.gds579
 PIN vccdgt_1p0.gds580
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 13.374 34.786 13.574 ;
 END
 END vccdgt_1p0.gds580
 PIN vccdgt_1p0.gds581
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.238 12.527 32.278 12.727 ;
 END
 END vccdgt_1p0.gds581
 PIN vccdgt_1p0.gds582
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.818 11.95 31.858 12.15 ;
 END
 END vccdgt_1p0.gds582
 PIN vccdgt_1p0.gds583
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.234 12.7505 31.29 12.9505 ;
 END
 END vccdgt_1p0.gds583
 PIN vccdgt_1p0.gds584
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.082 14.161 33.128 14.361 ;
 END
 END vccdgt_1p0.gds584
 PIN vccdgt_1p0.gds585
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.366 14.213 32.406 14.413 ;
 END
 END vccdgt_1p0.gds585
 PIN vccdgt_1p0.gds586
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.654 13.638 31.71 13.838 ;
 END
 END vccdgt_1p0.gds586
 PIN vccdgt_1p0.gds587
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.01 14.05 32.05 14.25 ;
 END
 END vccdgt_1p0.gds587
 PIN vccdgt_1p0.gds588
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.166 13.2825 35.226 13.4825 ;
 END
 END vccdgt_1p0.gds588
 PIN vccdgt_1p0.gds589
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.91 11.6505 34.95 11.8505 ;
 END
 END vccdgt_1p0.gds589
 PIN vccdgt_1p0.gds590
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.054 13.803 31.13 14.003 ;
 END
 END vccdgt_1p0.gds590
 PIN vccdgt_1p0.gds591
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.554 10.8945 30.61 11.0945 ;
 END
 END vccdgt_1p0.gds591
 PIN vccdgt_1p0.gds592
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.23 13.0715 34.286 13.2715 ;
 END
 END vccdgt_1p0.gds592
 PIN vccdgt_1p0.gds593
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.65 11.025 34.706 11.225 ;
 END
 END vccdgt_1p0.gds593
 PIN vccdgt_1p0.gds594
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.574 12.3155 32.634 12.5155 ;
 END
 END vccdgt_1p0.gds594
 PIN vccdgt_1p0.gds595
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.386 13.268 33.442 13.468 ;
 END
 END vccdgt_1p0.gds595
 PIN vccdgt_1p0.gds596
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.726 12.968 33.786 13.168 ;
 END
 END vccdgt_1p0.gds596
 PIN vccdgt_1p0.gds597
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 30.464 15.127 30.52 15.309 ;
 RECT 31.136 15.127 31.192 15.309 ;
 RECT 30.8 15.127 30.856 15.309 ;
 RECT 32.144 15.09 32.2 15.29 ;
 RECT 31.808 15.09 31.864 15.29 ;
 RECT 32.48 15.09 32.536 15.29 ;
 RECT 33.74 15.109 33.796 15.309 ;
 RECT 33.32 15.127 33.376 15.309 ;
 RECT 34.832 15.091 34.888 15.291 ;
 RECT 32.312 15.37 32.368 15.57 ;
 RECT 30.632 15.37 30.688 15.57 ;
 RECT 30.296 15.3035 30.352 15.5035 ;
 RECT 30.968 15.2705 31.024 15.4705 ;
 RECT 31.976 15.37 32.032 15.57 ;
 RECT 32.984 15.37 33.04 15.57 ;
 RECT 32.648 15.37 32.704 15.57 ;
 RECT 33.32 15.37 33.376 15.57 ;
 RECT 34.58 15.23 34.636 15.43 ;
 RECT 34.244 15.351 34.3 15.533 ;
 RECT 34.832 15.369 34.888 15.569 ;
 RECT 30.464 14.007 30.52 14.189 ;
 RECT 30.296 13.989 30.352 14.189 ;
 RECT 31.304 14.007 31.36 14.189 ;
 RECT 31.136 14.007 31.192 14.189 ;
 RECT 30.8 14.007 30.856 14.189 ;
 RECT 32.144 14.026 32.2 14.226 ;
 RECT 31.808 14.026 31.864 14.226 ;
 RECT 31.64 14.007 31.696 14.189 ;
 RECT 32.48 14.026 32.536 14.226 ;
 RECT 32.984 14.007 33.04 14.189 ;
 RECT 32.816 14.007 32.872 14.189 ;
 RECT 33.74 14.007 33.796 14.189 ;
 RECT 33.572 14.007 33.628 14.189 ;
 RECT 33.404 14.007 33.46 14.189 ;
 RECT 34.412 14.007 34.468 14.189 ;
 RECT 34.244 14.007 34.3 14.189 ;
 RECT 35.168 14.064 35.224 14.264 ;
 RECT 30.548 12.682 30.604 12.882 ;
 RECT 32.228 12.682 32.284 12.882 ;
 RECT 31.892 12.682 31.948 12.882 ;
 RECT 33.152 12.679 33.208 12.843 ;
 RECT 32.564 12.682 32.62 12.882 ;
 RECT 32.9 12.672 32.956 12.843 ;
 RECT 34.58 12.681 34.636 12.881 ;
 RECT 30.464 12.439 30.52 12.621 ;
 RECT 30.296 12.439 30.352 12.621 ;
 RECT 31.388 12.542 31.444 12.742 ;
 RECT 31.136 12.439 31.192 12.621 ;
 RECT 30.968 12.542 31.024 12.742 ;
 RECT 30.8 12.439 30.856 12.621 ;
 RECT 31.892 12.402 31.948 12.602 ;
 RECT 31.724 12.542 31.78 12.742 ;
 RECT 32.984 12.439 33.04 12.621 ;
 RECT 32.816 12.439 32.872 12.621 ;
 RECT 32.648 12.439 32.704 12.621 ;
 RECT 32.48 12.439 32.536 12.621 ;
 RECT 33.656 12.403 33.712 12.603 ;
 RECT 33.236 12.441 33.292 12.621 ;
 RECT 34.58 12.403 34.636 12.603 ;
 RECT 33.992 12.402 34.048 12.602 ;
 RECT 34.832 12.403 34.888 12.603 ;
 RECT 30.464 11.319 30.52 11.501 ;
 RECT 30.296 11.319 30.352 11.501 ;
 RECT 31.388 11.319 31.444 11.501 ;
 RECT 31.136 11.319 31.192 11.501 ;
 RECT 30.968 11.319 31.024 11.501 ;
 RECT 30.8 11.319 30.856 11.501 ;
 RECT 31.892 11.319 31.948 11.501 ;
 RECT 31.724 11.301 31.78 11.501 ;
 RECT 32.816 11.301 32.872 11.501 ;
 RECT 32.648 11.301 32.704 11.501 ;
 RECT 32.48 11.301 32.536 11.501 ;
 RECT 33.74 11.338 33.796 11.538 ;
 RECT 33.572 11.301 33.628 11.501 ;
 RECT 33.404 11.301 33.46 11.501 ;
 RECT 34.58 11.301 34.636 11.501 ;
 RECT 34.916 11.337 34.972 11.537 ;
 RECT 31.976 11.058 32.032 11.258 ;
 RECT 31.64 11.058 31.696 11.258 ;
 RECT 30.968 11.058 31.024 11.258 ;
 RECT 30.632 11.058 30.688 11.258 ;
 RECT 30.296 11.058 30.352 11.258 ;
 RECT 33.656 11.058 33.712 11.258 ;
 RECT 33.992 11.058 34.048 11.258 ;
 RECT 30.548 13.676 30.604 13.876 ;
 RECT 31.388 13.676 31.444 13.876 ;
 RECT 30.968 13.7925 31.024 13.9925 ;
 RECT 32.228 13.746 32.284 13.946 ;
 RECT 31.892 13.746 31.948 13.946 ;
 RECT 31.724 13.783 31.78 13.965 ;
 RECT 33.152 13.8845 33.208 14.0845 ;
 RECT 32.564 13.746 32.62 13.946 ;
 RECT 32.9 13.785 32.956 13.951 ;
 RECT 34.16 12.3615 34.216 12.5615 ;
 RECT 34.328 12.3615 34.384 12.5615 ;
 RECT 34.748 11.267 34.804 11.467 ;
 RECT 33.992 11.408 34.048 11.608 ;
 RECT 34.328 11.291 34.384 11.491 ;
 RECT 34.16 11.408 34.216 11.608 ;
 RECT 31.304 10.988 31.36 11.188 ;
 RECT 33.32 10.988 33.376 11.188 ;
 RECT 32.984 11.1275 33.04 11.3275 ;
 RECT 33.236 11.2685 33.292 11.4685 ;
 RECT 34.076 12.752 34.132 12.952 ;
 RECT 33.572 12.752 33.628 12.952 ;
 RECT 31.304 15.249 31.36 15.449 ;
 RECT 33.572 15.127 33.628 15.309 ;
 RECT 34.496 15.239 34.552 15.439 ;
 RECT 33.992 15.351 34.048 15.533 ;
 RECT 31.556 15.2025 31.612 15.4025 ;
 RECT 32.9 15.02 32.956 15.22 ;
 RECT 34.328 15.02 34.384 15.22 ;
 RECT 34.16 15.02 34.216 15.22 ;
 RECT 33.068 15.09 33.124 15.29 ;
 RECT 35.084 14.5165 35.14 14.7165 ;
 RECT 33.656 13.676 33.712 13.876 ;
 RECT 34.58 13.7265 34.636 13.9265 ;
 RECT 34.16 13.676 34.216 13.876 ;
 END
 END vccdgt_1p0.gds597
 PIN vccdgt_1p0.gds598
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.122 11.011 40.182 11.211 ;
 END
 END vccdgt_1p0.gds598
 PIN vccdgt_1p0.gds599
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.45 11.011 39.51 11.211 ;
 END
 END vccdgt_1p0.gds599
 PIN vccdgt_1p0.gds600
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.778 11.011 38.838 11.211 ;
 END
 END vccdgt_1p0.gds600
 PIN vccdgt_1p0.gds601
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.106 11.011 38.166 11.211 ;
 END
 END vccdgt_1p0.gds601
 PIN vccdgt_1p0.gds602
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.434 11.011 37.494 11.211 ;
 END
 END vccdgt_1p0.gds602
 PIN vccdgt_1p0.gds603
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.762 11.011 36.822 11.211 ;
 END
 END vccdgt_1p0.gds603
 PIN vccdgt_1p0.gds604
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.09 11.011 36.15 11.211 ;
 END
 END vccdgt_1p0.gds604
 PIN vccdgt_1p0.gds605
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.418 11.011 35.478 11.211 ;
 END
 END vccdgt_1p0.gds605
 PIN vccdgt_1p0.gds606
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.618 11.011 39.678 11.211 ;
 END
 END vccdgt_1p0.gds606
 PIN vccdgt_1p0.gds607
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.786 11.011 39.846 11.211 ;
 END
 END vccdgt_1p0.gds607
 PIN vccdgt_1p0.gds608
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.946 11.011 39.006 11.211 ;
 END
 END vccdgt_1p0.gds608
 PIN vccdgt_1p0.gds609
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.114 11.011 39.174 11.211 ;
 END
 END vccdgt_1p0.gds609
 PIN vccdgt_1p0.gds610
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.274 11.011 38.334 11.211 ;
 END
 END vccdgt_1p0.gds610
 PIN vccdgt_1p0.gds611
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.442 11.011 38.502 11.211 ;
 END
 END vccdgt_1p0.gds611
 PIN vccdgt_1p0.gds612
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.602 11.011 37.662 11.211 ;
 END
 END vccdgt_1p0.gds612
 PIN vccdgt_1p0.gds613
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.77 11.011 37.83 11.211 ;
 END
 END vccdgt_1p0.gds613
 PIN vccdgt_1p0.gds614
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.93 11.011 36.99 11.211 ;
 END
 END vccdgt_1p0.gds614
 PIN vccdgt_1p0.gds615
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.098 11.011 37.158 11.211 ;
 END
 END vccdgt_1p0.gds615
 PIN vccdgt_1p0.gds616
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.258 11.011 36.318 11.211 ;
 END
 END vccdgt_1p0.gds616
 PIN vccdgt_1p0.gds617
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.426 11.011 36.486 11.211 ;
 END
 END vccdgt_1p0.gds617
 PIN vccdgt_1p0.gds618
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.586 11.011 35.646 11.211 ;
 END
 END vccdgt_1p0.gds618
 PIN vccdgt_1p0.gds619
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.754 11.011 35.814 11.211 ;
 END
 END vccdgt_1p0.gds619
 PIN vccdgt_1p0.gds620
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.038 12.7505 40.078 12.9505 ;
 END
 END vccdgt_1p0.gds620
 PIN vccdgt_1p0.gds621
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.366 12.7505 39.406 12.9505 ;
 END
 END vccdgt_1p0.gds621
 PIN vccdgt_1p0.gds622
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.694 12.7505 38.734 12.9505 ;
 END
 END vccdgt_1p0.gds622
 PIN vccdgt_1p0.gds623
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.022 12.7505 38.062 12.9505 ;
 END
 END vccdgt_1p0.gds623
 PIN vccdgt_1p0.gds624
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.35 12.7505 37.39 12.9505 ;
 END
 END vccdgt_1p0.gds624
 PIN vccdgt_1p0.gds625
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.678 12.7505 36.718 12.9505 ;
 END
 END vccdgt_1p0.gds625
 PIN vccdgt_1p0.gds626
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.006 12.7505 36.046 12.9505 ;
 END
 END vccdgt_1p0.gds626
 PIN vccdgt_1p0.gds627
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.334 12.7505 35.374 12.9505 ;
 END
 END vccdgt_1p0.gds627
 PIN vccdgt_1p0.gds628
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.762 15.406 39.802 15.606 ;
 END
 END vccdgt_1p0.gds628
 PIN vccdgt_1p0.gds629
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.09 15.406 39.13 15.606 ;
 END
 END vccdgt_1p0.gds629
 PIN vccdgt_1p0.gds630
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.418 15.406 38.458 15.606 ;
 END
 END vccdgt_1p0.gds630
 PIN vccdgt_1p0.gds631
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.746 15.406 37.786 15.606 ;
 END
 END vccdgt_1p0.gds631
 PIN vccdgt_1p0.gds632
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.074 15.406 37.114 15.606 ;
 END
 END vccdgt_1p0.gds632
 PIN vccdgt_1p0.gds633
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.402 15.406 36.442 15.606 ;
 END
 END vccdgt_1p0.gds633
 PIN vccdgt_1p0.gds634
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.762 11.9905 39.802 12.1905 ;
 END
 END vccdgt_1p0.gds634
 PIN vccdgt_1p0.gds635
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.09 11.9905 39.13 12.1905 ;
 END
 END vccdgt_1p0.gds635
 PIN vccdgt_1p0.gds636
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.418 11.9905 38.458 12.1905 ;
 END
 END vccdgt_1p0.gds636
 PIN vccdgt_1p0.gds637
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.746 11.9905 37.786 12.1905 ;
 END
 END vccdgt_1p0.gds637
 PIN vccdgt_1p0.gds638
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.074 11.9905 37.114 12.1905 ;
 END
 END vccdgt_1p0.gds638
 PIN vccdgt_1p0.gds639
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.402 11.9905 36.442 12.1905 ;
 END
 END vccdgt_1p0.gds639
 PIN vccdgt_1p0.gds640
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.538 12.617 35.578 12.817 ;
 END
 END vccdgt_1p0.gds640
 PIN vccdgt_1p0.gds641
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.242 12.617 40.282 12.817 ;
 END
 END vccdgt_1p0.gds641
 PIN vccdgt_1p0.gds642
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.89 13.483 39.93 13.683 ;
 END
 END vccdgt_1p0.gds642
 PIN vccdgt_1p0.gds643
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.57 12.617 39.61 12.817 ;
 END
 END vccdgt_1p0.gds643
 PIN vccdgt_1p0.gds644
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.218 13.483 39.258 13.683 ;
 END
 END vccdgt_1p0.gds644
 PIN vccdgt_1p0.gds645
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.898 12.617 38.938 12.817 ;
 END
 END vccdgt_1p0.gds645
 PIN vccdgt_1p0.gds646
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.546 13.483 38.586 13.683 ;
 END
 END vccdgt_1p0.gds646
 PIN vccdgt_1p0.gds647
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.226 12.617 38.266 12.817 ;
 END
 END vccdgt_1p0.gds647
 PIN vccdgt_1p0.gds648
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.874 13.483 37.914 13.683 ;
 END
 END vccdgt_1p0.gds648
 PIN vccdgt_1p0.gds649
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.554 12.617 37.594 12.817 ;
 END
 END vccdgt_1p0.gds649
 PIN vccdgt_1p0.gds650
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.202 13.483 37.242 13.683 ;
 END
 END vccdgt_1p0.gds650
 PIN vccdgt_1p0.gds651
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.882 12.617 36.922 12.817 ;
 END
 END vccdgt_1p0.gds651
 PIN vccdgt_1p0.gds652
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.53 13.483 36.57 13.683 ;
 END
 END vccdgt_1p0.gds652
 PIN vccdgt_1p0.gds653
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.21 12.617 36.25 12.817 ;
 END
 END vccdgt_1p0.gds653
 PIN vccdgt_1p0.gds654
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.858 13.483 35.898 13.683 ;
 END
 END vccdgt_1p0.gds654
 PIN vccdgt_1p0.gds655
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.73 11.9905 35.77 12.1905 ;
 END
 END vccdgt_1p0.gds655
 PIN vccdgt_1p0.gds656
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.73 15.406 35.77 15.606 ;
 END
 END vccdgt_1p0.gds656
 PIN vccdgt_1p0.gds657
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 39.956 15.23 40.012 15.43 ;
 RECT 39.284 15.23 39.34 15.43 ;
 RECT 38.612 15.23 38.668 15.43 ;
 RECT 37.94 15.23 37.996 15.43 ;
 RECT 37.268 15.23 37.324 15.43 ;
 RECT 36.596 15.23 36.652 15.43 ;
 RECT 35.252 15.23 35.308 15.43 ;
 RECT 35.924 15.23 35.98 15.43 ;
 RECT 40.124 12.165 40.18 12.365 ;
 RECT 39.62 12.165 39.676 12.365 ;
 RECT 39.452 12.165 39.508 12.365 ;
 RECT 39.788 12.165 39.844 12.365 ;
 RECT 39.956 12.1635 40.012 12.3635 ;
 RECT 38.948 12.165 39.004 12.365 ;
 RECT 38.78 12.165 38.836 12.365 ;
 RECT 39.116 12.165 39.172 12.365 ;
 RECT 39.284 12.1635 39.34 12.3635 ;
 RECT 38.276 12.165 38.332 12.365 ;
 RECT 38.108 12.165 38.164 12.365 ;
 RECT 38.444 12.165 38.5 12.365 ;
 RECT 38.612 12.1635 38.668 12.3635 ;
 RECT 37.604 12.165 37.66 12.365 ;
 RECT 37.436 12.165 37.492 12.365 ;
 RECT 37.772 12.165 37.828 12.365 ;
 RECT 37.94 12.1635 37.996 12.3635 ;
 RECT 36.932 12.165 36.988 12.365 ;
 RECT 36.764 12.165 36.82 12.365 ;
 RECT 37.1 12.165 37.156 12.365 ;
 RECT 37.268 12.1635 37.324 12.3635 ;
 RECT 36.26 12.165 36.316 12.365 ;
 RECT 36.092 12.165 36.148 12.365 ;
 RECT 36.428 12.165 36.484 12.365 ;
 RECT 36.596 12.1635 36.652 12.3635 ;
 RECT 35.588 12.165 35.644 12.365 ;
 RECT 35.42 12.165 35.476 12.365 ;
 RECT 35.756 12.165 35.812 12.365 ;
 RECT 35.924 12.1635 35.98 12.3635 ;
 RECT 40.124 13.197 40.18 13.397 ;
 RECT 39.62 13.197 39.676 13.397 ;
 RECT 39.452 13.197 39.508 13.397 ;
 RECT 39.956 13.214 40.012 13.414 ;
 RECT 39.788 13.197 39.844 13.397 ;
 RECT 38.948 13.197 39.004 13.397 ;
 RECT 38.78 13.197 38.836 13.397 ;
 RECT 39.284 13.214 39.34 13.414 ;
 RECT 39.116 13.197 39.172 13.397 ;
 RECT 38.276 13.197 38.332 13.397 ;
 RECT 38.108 13.197 38.164 13.397 ;
 RECT 38.612 13.214 38.668 13.414 ;
 RECT 38.444 13.197 38.5 13.397 ;
 RECT 37.604 13.197 37.66 13.397 ;
 RECT 37.436 13.197 37.492 13.397 ;
 RECT 37.94 13.214 37.996 13.414 ;
 RECT 37.772 13.197 37.828 13.397 ;
 RECT 36.932 13.197 36.988 13.397 ;
 RECT 36.764 13.197 36.82 13.397 ;
 RECT 37.268 13.214 37.324 13.414 ;
 RECT 37.1 13.197 37.156 13.397 ;
 RECT 36.26 13.197 36.316 13.397 ;
 RECT 36.092 13.197 36.148 13.397 ;
 RECT 36.596 13.214 36.652 13.414 ;
 RECT 36.428 13.197 36.484 13.397 ;
 RECT 35.588 13.197 35.644 13.397 ;
 RECT 35.42 13.197 35.476 13.397 ;
 RECT 35.252 13.214 35.308 13.414 ;
 RECT 35.924 13.214 35.98 13.414 ;
 RECT 35.756 13.197 35.812 13.397 ;
 END
 END vccdgt_1p0.gds657
 PIN vccdgt_1p0.gds658
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.574 11.011 44.634 11.211 ;
 END
 END vccdgt_1p0.gds658
 PIN vccdgt_1p0.gds659
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.902 11.011 43.962 11.211 ;
 END
 END vccdgt_1p0.gds659
 PIN vccdgt_1p0.gds660
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.23 11.011 43.29 11.211 ;
 END
 END vccdgt_1p0.gds660
 PIN vccdgt_1p0.gds661
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.558 11.011 42.618 11.211 ;
 END
 END vccdgt_1p0.gds661
 PIN vccdgt_1p0.gds662
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.886 11.011 41.946 11.211 ;
 END
 END vccdgt_1p0.gds662
 PIN vccdgt_1p0.gds663
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.214 11.011 41.274 11.211 ;
 END
 END vccdgt_1p0.gds663
 PIN vccdgt_1p0.gds664
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.742 11.011 44.802 11.211 ;
 END
 END vccdgt_1p0.gds664
 PIN vccdgt_1p0.gds665
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.91 11.011 44.97 11.211 ;
 END
 END vccdgt_1p0.gds665
 PIN vccdgt_1p0.gds666
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.07 11.011 44.13 11.211 ;
 END
 END vccdgt_1p0.gds666
 PIN vccdgt_1p0.gds667
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.238 11.011 44.298 11.211 ;
 END
 END vccdgt_1p0.gds667
 PIN vccdgt_1p0.gds668
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.398 11.011 43.458 11.211 ;
 END
 END vccdgt_1p0.gds668
 PIN vccdgt_1p0.gds669
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.566 11.011 43.626 11.211 ;
 END
 END vccdgt_1p0.gds669
 PIN vccdgt_1p0.gds670
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.726 11.011 42.786 11.211 ;
 END
 END vccdgt_1p0.gds670
 PIN vccdgt_1p0.gds671
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.894 11.011 42.954 11.211 ;
 END
 END vccdgt_1p0.gds671
 PIN vccdgt_1p0.gds672
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.054 11.011 42.114 11.211 ;
 END
 END vccdgt_1p0.gds672
 PIN vccdgt_1p0.gds673
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.222 11.011 42.282 11.211 ;
 END
 END vccdgt_1p0.gds673
 PIN vccdgt_1p0.gds674
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.382 11.011 41.442 11.211 ;
 END
 END vccdgt_1p0.gds674
 PIN vccdgt_1p0.gds675
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.55 11.011 41.61 11.211 ;
 END
 END vccdgt_1p0.gds675
 PIN vccdgt_1p0.gds676
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.29 11.011 40.35 11.211 ;
 END
 END vccdgt_1p0.gds676
 PIN vccdgt_1p0.gds677
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.458 11.011 40.518 11.211 ;
 END
 END vccdgt_1p0.gds677
 PIN vccdgt_1p0.gds678
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.162 12.7505 45.202 12.9505 ;
 END
 END vccdgt_1p0.gds678
 PIN vccdgt_1p0.gds679
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.49 12.7505 44.53 12.9505 ;
 END
 END vccdgt_1p0.gds679
 PIN vccdgt_1p0.gds680
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.818 12.7505 43.858 12.9505 ;
 END
 END vccdgt_1p0.gds680
 PIN vccdgt_1p0.gds681
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.146 12.7505 43.186 12.9505 ;
 END
 END vccdgt_1p0.gds681
 PIN vccdgt_1p0.gds682
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.474 12.7505 42.514 12.9505 ;
 END
 END vccdgt_1p0.gds682
 PIN vccdgt_1p0.gds683
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.802 12.7505 41.842 12.9505 ;
 END
 END vccdgt_1p0.gds683
 PIN vccdgt_1p0.gds684
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.13 12.7505 41.17 12.9505 ;
 END
 END vccdgt_1p0.gds684
 PIN vccdgt_1p0.gds685
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.562 13.309 40.602 13.509 ;
 END
 END vccdgt_1p0.gds685
 PIN vccdgt_1p0.gds686
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.886 15.406 44.926 15.606 ;
 END
 END vccdgt_1p0.gds686
 PIN vccdgt_1p0.gds687
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.214 15.406 44.254 15.606 ;
 END
 END vccdgt_1p0.gds687
 PIN vccdgt_1p0.gds688
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.542 15.406 43.582 15.606 ;
 END
 END vccdgt_1p0.gds688
 PIN vccdgt_1p0.gds689
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.87 15.406 42.91 15.606 ;
 END
 END vccdgt_1p0.gds689
 PIN vccdgt_1p0.gds690
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.198 15.406 42.238 15.606 ;
 END
 END vccdgt_1p0.gds690
 PIN vccdgt_1p0.gds691
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.886 11.9905 44.926 12.1905 ;
 END
 END vccdgt_1p0.gds691
 PIN vccdgt_1p0.gds692
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.214 11.9905 44.254 12.1905 ;
 END
 END vccdgt_1p0.gds692
 PIN vccdgt_1p0.gds693
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.542 11.9905 43.582 12.1905 ;
 END
 END vccdgt_1p0.gds693
 PIN vccdgt_1p0.gds694
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.87 11.9905 42.91 12.1905 ;
 END
 END vccdgt_1p0.gds694
 PIN vccdgt_1p0.gds695
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.198 11.9905 42.238 12.1905 ;
 END
 END vccdgt_1p0.gds695
 PIN vccdgt_1p0.gds696
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.526 11.9905 41.566 12.1905 ;
 END
 END vccdgt_1p0.gds696
 PIN vccdgt_1p0.gds697
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.434 11.9905 40.474 12.1905 ;
 END
 END vccdgt_1p0.gds697
 PIN vccdgt_1p0.gds698
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.014 13.483 45.054 13.683 ;
 END
 END vccdgt_1p0.gds698
 PIN vccdgt_1p0.gds699
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.694 12.617 44.734 12.817 ;
 END
 END vccdgt_1p0.gds699
 PIN vccdgt_1p0.gds700
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.342 13.483 44.382 13.683 ;
 END
 END vccdgt_1p0.gds700
 PIN vccdgt_1p0.gds701
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.022 12.617 44.062 12.817 ;
 END
 END vccdgt_1p0.gds701
 PIN vccdgt_1p0.gds702
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.67 13.483 43.71 13.683 ;
 END
 END vccdgt_1p0.gds702
 PIN vccdgt_1p0.gds703
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.35 12.617 43.39 12.817 ;
 END
 END vccdgt_1p0.gds703
 PIN vccdgt_1p0.gds704
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.998 13.483 43.038 13.683 ;
 END
 END vccdgt_1p0.gds704
 PIN vccdgt_1p0.gds705
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.678 12.617 42.718 12.817 ;
 END
 END vccdgt_1p0.gds705
 PIN vccdgt_1p0.gds706
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.326 13.483 42.366 13.683 ;
 END
 END vccdgt_1p0.gds706
 PIN vccdgt_1p0.gds707
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.006 12.617 42.046 12.817 ;
 END
 END vccdgt_1p0.gds707
 PIN vccdgt_1p0.gds708
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.654 13.483 41.694 13.683 ;
 END
 END vccdgt_1p0.gds708
 PIN vccdgt_1p0.gds709
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.334 12.617 41.374 12.817 ;
 END
 END vccdgt_1p0.gds709
 PIN vccdgt_1p0.gds710
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.982 13.4245 41.022 13.6245 ;
 END
 END vccdgt_1p0.gds710
 PIN vccdgt_1p0.gds711
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.71 13.0135 40.75 13.2135 ;
 END
 END vccdgt_1p0.gds711
 PIN vccdgt_1p0.gds712
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.526 15.406 41.566 15.606 ;
 END
 END vccdgt_1p0.gds712
 PIN vccdgt_1p0.gds713
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.434 15.406 40.474 15.606 ;
 END
 END vccdgt_1p0.gds713
 PIN vccdgt_1p0.gds714
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 45.08 15.23 45.136 15.43 ;
 RECT 44.408 15.23 44.464 15.43 ;
 RECT 43.736 15.23 43.792 15.43 ;
 RECT 43.064 15.23 43.12 15.43 ;
 RECT 42.392 15.23 42.448 15.43 ;
 RECT 41.048 15.23 41.104 15.43 ;
 RECT 41.72 15.23 41.776 15.43 ;
 RECT 40.628 15.23 40.684 15.43 ;
 RECT 44.744 12.165 44.8 12.365 ;
 RECT 44.576 12.165 44.632 12.365 ;
 RECT 44.912 12.165 44.968 12.365 ;
 RECT 45.08 12.1635 45.136 12.3635 ;
 RECT 44.072 12.165 44.128 12.365 ;
 RECT 43.904 12.165 43.96 12.365 ;
 RECT 44.24 12.165 44.296 12.365 ;
 RECT 44.408 12.1635 44.464 12.3635 ;
 RECT 43.4 12.165 43.456 12.365 ;
 RECT 43.232 12.165 43.288 12.365 ;
 RECT 43.568 12.165 43.624 12.365 ;
 RECT 43.736 12.1635 43.792 12.3635 ;
 RECT 42.728 12.165 42.784 12.365 ;
 RECT 42.56 12.165 42.616 12.365 ;
 RECT 42.896 12.165 42.952 12.365 ;
 RECT 43.064 12.1635 43.12 12.3635 ;
 RECT 42.056 12.165 42.112 12.365 ;
 RECT 41.888 12.165 41.944 12.365 ;
 RECT 42.224 12.165 42.28 12.365 ;
 RECT 42.392 12.1635 42.448 12.3635 ;
 RECT 41.384 12.165 41.44 12.365 ;
 RECT 41.216 12.165 41.272 12.365 ;
 RECT 41.552 12.165 41.608 12.365 ;
 RECT 41.72 12.1635 41.776 12.3635 ;
 RECT 40.46 12.165 40.516 12.365 ;
 RECT 40.628 12.1635 40.684 12.3635 ;
 RECT 40.292 12.165 40.348 12.365 ;
 RECT 40.88 13.659 40.936 13.859 ;
 RECT 40.964 13.095 41.02 13.295 ;
 RECT 40.712 13.2495 40.768 13.4495 ;
 RECT 44.744 13.197 44.8 13.397 ;
 RECT 44.576 13.197 44.632 13.397 ;
 RECT 45.08 13.214 45.136 13.414 ;
 RECT 44.912 13.197 44.968 13.397 ;
 RECT 44.072 13.197 44.128 13.397 ;
 RECT 43.904 13.197 43.96 13.397 ;
 RECT 44.408 13.214 44.464 13.414 ;
 RECT 44.24 13.197 44.296 13.397 ;
 RECT 43.4 13.197 43.456 13.397 ;
 RECT 43.232 13.197 43.288 13.397 ;
 RECT 43.736 13.214 43.792 13.414 ;
 RECT 43.568 13.197 43.624 13.397 ;
 RECT 42.728 13.197 42.784 13.397 ;
 RECT 42.56 13.197 42.616 13.397 ;
 RECT 43.064 13.214 43.12 13.414 ;
 RECT 42.896 13.197 42.952 13.397 ;
 RECT 42.056 13.197 42.112 13.397 ;
 RECT 41.888 13.197 41.944 13.397 ;
 RECT 42.392 13.214 42.448 13.414 ;
 RECT 42.224 13.197 42.28 13.397 ;
 RECT 41.384 13.197 41.44 13.397 ;
 RECT 41.216 13.197 41.272 13.397 ;
 RECT 41.048 13.214 41.104 13.414 ;
 RECT 41.72 13.214 41.776 13.414 ;
 RECT 41.552 13.197 41.608 13.397 ;
 RECT 40.628 13.214 40.684 13.414 ;
 RECT 40.46 13.197 40.516 13.397 ;
 RECT 40.292 13.197 40.348 13.397 ;
 END
 END vccdgt_1p0.gds714
 PIN vccdgt_1p0.gds715
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.918 11.011 45.978 11.211 ;
 END
 END vccdgt_1p0.gds715
 PIN vccdgt_1p0.gds716
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.246 11.011 45.306 11.211 ;
 END
 END vccdgt_1p0.gds716
 PIN vccdgt_1p0.gds717
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.526 15.003 47.582 15.203 ;
 END
 END vccdgt_1p0.gds717
 PIN vccdgt_1p0.gds718
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.446 10.662 47.502 10.862 ;
 END
 END vccdgt_1p0.gds718
 PIN vccdgt_1p0.gds719
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.97 14.062 50.03 14.262 ;
 END
 END vccdgt_1p0.gds719
 PIN vccdgt_1p0.gds720
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.086 11.011 46.146 11.211 ;
 END
 END vccdgt_1p0.gds720
 PIN vccdgt_1p0.gds721
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.254 11.011 46.314 11.211 ;
 END
 END vccdgt_1p0.gds721
 PIN vccdgt_1p0.gds722
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.414 11.011 45.474 11.211 ;
 END
 END vccdgt_1p0.gds722
 PIN vccdgt_1p0.gds723
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.582 11.011 45.642 11.211 ;
 END
 END vccdgt_1p0.gds723
 PIN vccdgt_1p0.gds724
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.358 13.309 46.398 13.509 ;
 END
 END vccdgt_1p0.gds724
 PIN vccdgt_1p0.gds725
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.834 12.7505 45.874 12.9505 ;
 END
 END vccdgt_1p0.gds725
 PIN vccdgt_1p0.gds726
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.558 15.406 45.598 15.606 ;
 END
 END vccdgt_1p0.gds726
 PIN vccdgt_1p0.gds727
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.23 11.9905 46.27 12.1905 ;
 END
 END vccdgt_1p0.gds727
 PIN vccdgt_1p0.gds728
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.558 11.9905 45.598 12.1905 ;
 END
 END vccdgt_1p0.gds728
 PIN vccdgt_1p0.gds729
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.038 12.617 46.078 12.817 ;
 END
 END vccdgt_1p0.gds729
 PIN vccdgt_1p0.gds730
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.686 13.483 45.726 13.683 ;
 END
 END vccdgt_1p0.gds730
 PIN vccdgt_1p0.gds731
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.366 12.617 45.406 12.817 ;
 END
 END vccdgt_1p0.gds731
 PIN vccdgt_1p0.gds732
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.606 10.8945 47.662 11.0945 ;
 END
 END vccdgt_1p0.gds732
 PIN vccdgt_1p0.gds733
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.026 11.224 47.082 11.424 ;
 END
 END vccdgt_1p0.gds733
 PIN vccdgt_1p0.gds734
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.418 14.213 49.458 14.413 ;
 END
 END vccdgt_1p0.gds734
 PIN vccdgt_1p0.gds735
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.706 13.638 48.762 13.838 ;
 END
 END vccdgt_1p0.gds735
 PIN vccdgt_1p0.gds736
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.026 14.7305 47.082 14.9305 ;
 END
 END vccdgt_1p0.gds736
 PIN vccdgt_1p0.gds737
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.266 13.189 47.342 13.389 ;
 END
 END vccdgt_1p0.gds737
 PIN vccdgt_1p0.gds738
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.106 13.803 48.182 14.003 ;
 END
 END vccdgt_1p0.gds738
 PIN vccdgt_1p0.gds739
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.23 15.406 46.27 15.606 ;
 END
 END vccdgt_1p0.gds739
 PIN vccdgt_1p0.gds740
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.29 12.527 49.33 12.727 ;
 END
 END vccdgt_1p0.gds740
 PIN vccdgt_1p0.gds741
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.87 11.95 48.91 12.15 ;
 END
 END vccdgt_1p0.gds741
 PIN vccdgt_1p0.gds742
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.286 12.7505 48.342 12.9505 ;
 END
 END vccdgt_1p0.gds742
 PIN vccdgt_1p0.gds743
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.626 12.3155 49.686 12.5155 ;
 END
 END vccdgt_1p0.gds743
 PIN vccdgt_1p0.gds744
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.062 14.05 49.102 14.25 ;
 END
 END vccdgt_1p0.gds744
 PIN vccdgt_1p0.gds745
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.134 14.161 50.18 14.361 ;
 END
 END vccdgt_1p0.gds745
 PIN vccdgt_1p0.gds746
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.782 10.478 46.822 10.678 ;
 END
 END vccdgt_1p0.gds746
 PIN vccdgt_1p0.gds747
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.506 13.446 46.566 13.646 ;
 END
 END vccdgt_1p0.gds747
 PIN vccdgt_1p0.gds748
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 46.844 15.091 46.9 15.291 ;
 RECT 47.18 15.127 47.236 15.309 ;
 RECT 47.516 15.127 47.572 15.309 ;
 RECT 48.188 15.127 48.244 15.309 ;
 RECT 47.852 15.127 47.908 15.309 ;
 RECT 49.196 15.09 49.252 15.29 ;
 RECT 48.86 15.09 48.916 15.29 ;
 RECT 49.532 15.09 49.588 15.29 ;
 RECT 49.364 15.37 49.42 15.57 ;
 RECT 46.844 15.37 46.9 15.57 ;
 RECT 47.684 15.37 47.74 15.57 ;
 RECT 47.348 15.3035 47.404 15.5035 ;
 RECT 47.012 15.4105 47.068 15.6105 ;
 RECT 48.02 15.2705 48.076 15.4705 ;
 RECT 49.028 15.37 49.084 15.57 ;
 RECT 50.036 15.37 50.092 15.57 ;
 RECT 49.7 15.37 49.756 15.57 ;
 RECT 46.424 15.23 46.48 15.43 ;
 RECT 45.752 15.23 45.808 15.43 ;
 RECT 47.516 14.007 47.572 14.189 ;
 RECT 47.348 13.989 47.404 14.189 ;
 RECT 48.356 14.007 48.412 14.189 ;
 RECT 48.188 14.007 48.244 14.189 ;
 RECT 47.852 14.007 47.908 14.189 ;
 RECT 49.196 14.026 49.252 14.226 ;
 RECT 48.86 14.026 48.916 14.226 ;
 RECT 48.692 14.007 48.748 14.189 ;
 RECT 49.532 14.026 49.588 14.226 ;
 RECT 50.036 14.007 50.092 14.189 ;
 RECT 49.868 14.007 49.924 14.189 ;
 RECT 47.6 12.682 47.656 12.882 ;
 RECT 47.18 12.682 47.236 12.882 ;
 RECT 49.28 12.682 49.336 12.882 ;
 RECT 48.944 12.682 49 12.882 ;
 RECT 50.204 12.679 50.26 12.843 ;
 RECT 49.616 12.682 49.672 12.882 ;
 RECT 49.952 12.672 50.008 12.843 ;
 RECT 46.76 12.403 46.816 12.603 ;
 RECT 47.516 12.439 47.572 12.621 ;
 RECT 47.348 12.439 47.404 12.621 ;
 RECT 47.18 12.439 47.236 12.621 ;
 RECT 48.44 12.542 48.496 12.742 ;
 RECT 48.188 12.439 48.244 12.621 ;
 RECT 48.02 12.542 48.076 12.742 ;
 RECT 47.852 12.439 47.908 12.621 ;
 RECT 48.944 12.402 49 12.602 ;
 RECT 48.776 12.542 48.832 12.742 ;
 RECT 50.036 12.439 50.092 12.621 ;
 RECT 49.868 12.439 49.924 12.621 ;
 RECT 49.7 12.439 49.756 12.621 ;
 RECT 49.532 12.439 49.588 12.621 ;
 RECT 46.76 11.337 46.816 11.537 ;
 RECT 47.18 11.319 47.236 11.501 ;
 RECT 47.516 11.319 47.572 11.501 ;
 RECT 47.348 11.319 47.404 11.501 ;
 RECT 48.44 11.319 48.496 11.501 ;
 RECT 48.188 11.319 48.244 11.501 ;
 RECT 48.02 11.319 48.076 11.501 ;
 RECT 47.852 11.319 47.908 11.501 ;
 RECT 48.944 11.319 49 11.501 ;
 RECT 48.776 11.301 48.832 11.501 ;
 RECT 49.868 11.301 49.924 11.501 ;
 RECT 49.7 11.301 49.756 11.501 ;
 RECT 49.532 11.301 49.588 11.501 ;
 RECT 49.028 11.058 49.084 11.258 ;
 RECT 48.692 11.058 48.748 11.258 ;
 RECT 47.012 11.058 47.068 11.258 ;
 RECT 48.02 11.058 48.076 11.258 ;
 RECT 47.684 11.058 47.74 11.258 ;
 RECT 47.348 11.058 47.404 11.258 ;
 RECT 46.76 11.059 46.816 11.259 ;
 RECT 47.6 13.676 47.656 13.876 ;
 RECT 47.18 13.886 47.236 14.086 ;
 RECT 48.44 13.676 48.496 13.876 ;
 RECT 48.02 13.7925 48.076 13.9925 ;
 RECT 49.28 13.746 49.336 13.946 ;
 RECT 48.944 13.746 49 13.946 ;
 RECT 48.776 13.783 48.832 13.965 ;
 RECT 50.204 13.8845 50.26 14.0845 ;
 RECT 49.616 13.746 49.672 13.946 ;
 RECT 49.952 13.785 50.008 13.951 ;
 RECT 48.356 10.988 48.412 11.188 ;
 RECT 47.012 13.634 47.068 13.834 ;
 RECT 46.676 14.1515 46.732 14.3515 ;
 RECT 50.036 11.1275 50.092 11.3275 ;
 RECT 48.356 15.249 48.412 15.449 ;
 RECT 48.608 15.2025 48.664 15.4025 ;
 RECT 49.952 15.02 50.008 15.22 ;
 RECT 50.12 15.09 50.176 15.29 ;
 RECT 46.088 12.165 46.144 12.365 ;
 RECT 45.92 12.165 45.976 12.365 ;
 RECT 46.256 12.165 46.312 12.365 ;
 RECT 46.424 12.1635 46.48 12.3635 ;
 RECT 45.416 12.165 45.472 12.365 ;
 RECT 45.248 12.165 45.304 12.365 ;
 RECT 45.584 12.165 45.64 12.365 ;
 RECT 45.752 12.1635 45.808 12.3635 ;
 RECT 46.088 13.197 46.144 13.397 ;
 RECT 45.92 13.197 45.976 13.397 ;
 RECT 46.424 13.214 46.48 13.414 ;
 RECT 46.256 13.197 46.312 13.397 ;
 RECT 45.416 13.197 45.472 13.397 ;
 RECT 45.248 13.197 45.304 13.397 ;
 RECT 45.752 13.214 45.808 13.414 ;
 RECT 45.584 13.197 45.64 13.397 ;
 END
 END vccdgt_1p0.gds748
 PIN vccdgt_1p0.gds749
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.158 11.011 55.218 11.211 ;
 END
 END vccdgt_1p0.gds749
 PIN vccdgt_1p0.gds750
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.486 11.011 54.546 11.211 ;
 END
 END vccdgt_1p0.gds750
 PIN vccdgt_1p0.gds751
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.814 11.011 53.874 11.211 ;
 END
 END vccdgt_1p0.gds751
 PIN vccdgt_1p0.gds752
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.142 11.011 53.202 11.211 ;
 END
 END vccdgt_1p0.gds752
 PIN vccdgt_1p0.gds753
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.47 11.011 52.53 11.211 ;
 END
 END vccdgt_1p0.gds753
 PIN vccdgt_1p0.gds754
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.074 12.7505 55.114 12.9505 ;
 END
 END vccdgt_1p0.gds754
 PIN vccdgt_1p0.gds755
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.402 12.7505 54.442 12.9505 ;
 END
 END vccdgt_1p0.gds755
 PIN vccdgt_1p0.gds756
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.73 12.7505 53.77 12.9505 ;
 END
 END vccdgt_1p0.gds756
 PIN vccdgt_1p0.gds757
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.122 13.1425 51.178 13.3425 ;
 END
 END vccdgt_1p0.gds757
 PIN vccdgt_1p0.gds758
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.942 12.5175 50.998 12.7175 ;
 END
 END vccdgt_1p0.gds758
 PIN vccdgt_1p0.gds759
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.654 11.011 54.714 11.211 ;
 END
 END vccdgt_1p0.gds759
 PIN vccdgt_1p0.gds760
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.822 11.011 54.882 11.211 ;
 END
 END vccdgt_1p0.gds760
 PIN vccdgt_1p0.gds761
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.982 11.011 54.042 11.211 ;
 END
 END vccdgt_1p0.gds761
 PIN vccdgt_1p0.gds762
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.15 11.011 54.21 11.211 ;
 END
 END vccdgt_1p0.gds762
 PIN vccdgt_1p0.gds763
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.31 11.011 53.37 11.211 ;
 END
 END vccdgt_1p0.gds763
 PIN vccdgt_1p0.gds764
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.478 11.011 53.538 11.211 ;
 END
 END vccdgt_1p0.gds764
 PIN vccdgt_1p0.gds765
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.638 11.011 52.698 11.211 ;
 END
 END vccdgt_1p0.gds765
 PIN vccdgt_1p0.gds766
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.806 11.011 52.866 11.211 ;
 END
 END vccdgt_1p0.gds766
 PIN vccdgt_1p0.gds767
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 10.502 50.674 10.702 ;
 END
 END vccdgt_1p0.gds767
 PIN vccdgt_1p0.gds768
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.058 12.7505 53.098 12.9505 ;
 END
 END vccdgt_1p0.gds768
 PIN vccdgt_1p0.gds769
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.386 12.7505 52.426 12.9505 ;
 END
 END vccdgt_1p0.gds769
 PIN vccdgt_1p0.gds770
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.798 15.406 54.838 15.606 ;
 END
 END vccdgt_1p0.gds770
 PIN vccdgt_1p0.gds771
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.126 15.406 54.166 15.606 ;
 END
 END vccdgt_1p0.gds771
 PIN vccdgt_1p0.gds772
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.454 15.406 53.494 15.606 ;
 END
 END vccdgt_1p0.gds772
 PIN vccdgt_1p0.gds773
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.438 13.268 50.494 13.468 ;
 END
 END vccdgt_1p0.gds773
 PIN vccdgt_1p0.gds774
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.442 13.2505 51.518 13.4505 ;
 END
 END vccdgt_1p0.gds774
 PIN vccdgt_1p0.gds775
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.778 12.968 50.838 13.168 ;
 END
 END vccdgt_1p0.gds775
 PIN vccdgt_1p0.gds776
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.59 12.617 52.63 12.817 ;
 END
 END vccdgt_1p0.gds776
 PIN vccdgt_1p0.gds777
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.278 12.617 55.318 12.817 ;
 END
 END vccdgt_1p0.gds777
 PIN vccdgt_1p0.gds778
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.926 13.483 54.966 13.683 ;
 END
 END vccdgt_1p0.gds778
 PIN vccdgt_1p0.gds779
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.606 12.617 54.646 12.817 ;
 END
 END vccdgt_1p0.gds779
 PIN vccdgt_1p0.gds780
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.254 13.483 54.294 13.683 ;
 END
 END vccdgt_1p0.gds780
 PIN vccdgt_1p0.gds781
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.798 11.9905 54.838 12.1905 ;
 END
 END vccdgt_1p0.gds781
 PIN vccdgt_1p0.gds782
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.934 12.617 53.974 12.817 ;
 END
 END vccdgt_1p0.gds782
 PIN vccdgt_1p0.gds783
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.582 13.483 53.622 13.683 ;
 END
 END vccdgt_1p0.gds783
 PIN vccdgt_1p0.gds784
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.126 11.9905 54.166 12.1905 ;
 END
 END vccdgt_1p0.gds784
 PIN vccdgt_1p0.gds785
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 13.374 51.838 13.574 ;
 END
 END vccdgt_1p0.gds785
 PIN vccdgt_1p0.gds786
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.962 11.6505 52.002 11.8505 ;
 END
 END vccdgt_1p0.gds786
 PIN vccdgt_1p0.gds787
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.702 11.025 51.758 11.225 ;
 END
 END vccdgt_1p0.gds787
 PIN vccdgt_1p0.gds788
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.262 12.617 53.302 12.817 ;
 END
 END vccdgt_1p0.gds788
 PIN vccdgt_1p0.gds789
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.91 13.483 52.95 13.683 ;
 END
 END vccdgt_1p0.gds789
 PIN vccdgt_1p0.gds790
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.454 11.9905 53.494 12.1905 ;
 END
 END vccdgt_1p0.gds790
 PIN vccdgt_1p0.gds791
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.782 11.9905 52.822 12.1905 ;
 END
 END vccdgt_1p0.gds791
 PIN vccdgt_1p0.gds792
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.218 13.2825 52.278 13.4825 ;
 END
 END vccdgt_1p0.gds792
 PIN vccdgt_1p0.gds793
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.282 13.0715 51.338 13.2715 ;
 END
 END vccdgt_1p0.gds793
 PIN vccdgt_1p0.gds794
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.782 15.406 52.822 15.606 ;
 END
 END vccdgt_1p0.gds794
 PIN vccdgt_1p0.gds795
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 50.792 15.109 50.848 15.309 ;
 RECT 50.372 15.127 50.428 15.309 ;
 RECT 51.884 15.091 51.94 15.291 ;
 RECT 54.992 15.23 55.048 15.43 ;
 RECT 54.32 15.23 54.376 15.43 ;
 RECT 50.372 15.37 50.428 15.57 ;
 RECT 51.632 15.23 51.688 15.43 ;
 RECT 51.296 15.351 51.352 15.533 ;
 RECT 51.884 15.369 51.94 15.569 ;
 RECT 53.648 15.23 53.704 15.43 ;
 RECT 52.304 15.23 52.36 15.43 ;
 RECT 52.976 15.23 53.032 15.43 ;
 RECT 50.792 14.007 50.848 14.189 ;
 RECT 50.624 14.007 50.68 14.189 ;
 RECT 50.456 14.007 50.512 14.189 ;
 RECT 51.464 14.007 51.52 14.189 ;
 RECT 51.296 14.007 51.352 14.189 ;
 RECT 52.22 14.064 52.276 14.264 ;
 RECT 51.632 12.681 51.688 12.881 ;
 RECT 50.708 12.403 50.764 12.603 ;
 RECT 50.288 12.441 50.344 12.621 ;
 RECT 51.632 12.403 51.688 12.603 ;
 RECT 51.044 12.402 51.1 12.602 ;
 RECT 51.884 12.403 51.94 12.603 ;
 RECT 50.792 11.338 50.848 11.538 ;
 RECT 50.624 11.301 50.68 11.501 ;
 RECT 50.456 11.301 50.512 11.501 ;
 RECT 51.632 11.301 51.688 11.501 ;
 RECT 51.968 11.337 52.024 11.537 ;
 RECT 50.708 11.058 50.764 11.258 ;
 RECT 51.044 11.058 51.1 11.258 ;
 RECT 51.212 12.3615 51.268 12.5615 ;
 RECT 51.38 12.3615 51.436 12.5615 ;
 RECT 51.044 11.408 51.1 11.608 ;
 RECT 51.38 11.291 51.436 11.491 ;
 RECT 51.212 11.408 51.268 11.608 ;
 RECT 51.128 12.752 51.184 12.952 ;
 RECT 50.624 12.752 50.68 12.952 ;
 RECT 50.372 10.988 50.428 11.188 ;
 RECT 50.288 11.2685 50.344 11.4685 ;
 RECT 50.708 13.676 50.764 13.876 ;
 RECT 51.632 13.7265 51.688 13.9265 ;
 RECT 51.212 13.676 51.268 13.876 ;
 RECT 51.8 11.267 51.856 11.467 ;
 RECT 55.16 12.165 55.216 12.365 ;
 RECT 54.656 12.165 54.712 12.365 ;
 RECT 54.488 12.165 54.544 12.365 ;
 RECT 54.824 12.165 54.88 12.365 ;
 RECT 54.992 12.1635 55.048 12.3635 ;
 RECT 53.984 12.165 54.04 12.365 ;
 RECT 53.816 12.165 53.872 12.365 ;
 RECT 54.152 12.165 54.208 12.365 ;
 RECT 54.32 12.1635 54.376 12.3635 ;
 RECT 53.312 12.165 53.368 12.365 ;
 RECT 53.144 12.165 53.2 12.365 ;
 RECT 53.48 12.165 53.536 12.365 ;
 RECT 53.648 12.1635 53.704 12.3635 ;
 RECT 52.64 12.165 52.696 12.365 ;
 RECT 52.472 12.165 52.528 12.365 ;
 RECT 52.808 12.165 52.864 12.365 ;
 RECT 52.976 12.1635 53.032 12.3635 ;
 RECT 52.136 14.5165 52.192 14.7165 ;
 RECT 50.624 15.127 50.68 15.309 ;
 RECT 51.548 15.239 51.604 15.439 ;
 RECT 51.044 15.351 51.1 15.533 ;
 RECT 51.38 15.02 51.436 15.22 ;
 RECT 51.212 15.02 51.268 15.22 ;
 RECT 55.16 13.197 55.216 13.397 ;
 RECT 54.656 13.197 54.712 13.397 ;
 RECT 54.488 13.197 54.544 13.397 ;
 RECT 54.992 13.214 55.048 13.414 ;
 RECT 54.824 13.197 54.88 13.397 ;
 RECT 53.984 13.197 54.04 13.397 ;
 RECT 53.816 13.197 53.872 13.397 ;
 RECT 54.32 13.214 54.376 13.414 ;
 RECT 54.152 13.197 54.208 13.397 ;
 RECT 53.312 13.197 53.368 13.397 ;
 RECT 53.144 13.197 53.2 13.397 ;
 RECT 53.648 13.214 53.704 13.414 ;
 RECT 53.48 13.197 53.536 13.397 ;
 RECT 52.64 13.197 52.696 13.397 ;
 RECT 52.472 13.197 52.528 13.397 ;
 RECT 52.304 13.214 52.36 13.414 ;
 RECT 52.976 13.214 53.032 13.414 ;
 RECT 52.808 13.197 52.864 13.397 ;
 END
 END vccdgt_1p0.gds795
 PIN vccdgt_1p0.gds796
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.61 11.011 59.67 11.211 ;
 END
 END vccdgt_1p0.gds796
 PIN vccdgt_1p0.gds797
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.938 11.011 58.998 11.211 ;
 END
 END vccdgt_1p0.gds797
 PIN vccdgt_1p0.gds798
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.266 11.011 58.326 11.211 ;
 END
 END vccdgt_1p0.gds798
 PIN vccdgt_1p0.gds799
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.174 11.011 57.234 11.211 ;
 END
 END vccdgt_1p0.gds799
 PIN vccdgt_1p0.gds800
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.502 11.011 56.562 11.211 ;
 END
 END vccdgt_1p0.gds800
 PIN vccdgt_1p0.gds801
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.83 11.011 55.89 11.211 ;
 END
 END vccdgt_1p0.gds801
 PIN vccdgt_1p0.gds802
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.614 13.309 57.654 13.509 ;
 END
 END vccdgt_1p0.gds802
 PIN vccdgt_1p0.gds803
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.198 12.7505 60.238 12.9505 ;
 END
 END vccdgt_1p0.gds803
 PIN vccdgt_1p0.gds804
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.526 12.7505 59.566 12.9505 ;
 END
 END vccdgt_1p0.gds804
 PIN vccdgt_1p0.gds805
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.854 12.7505 58.894 12.9505 ;
 END
 END vccdgt_1p0.gds805
 PIN vccdgt_1p0.gds806
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.182 12.7505 58.222 12.9505 ;
 END
 END vccdgt_1p0.gds806
 PIN vccdgt_1p0.gds807
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.09 12.7505 57.13 12.9505 ;
 END
 END vccdgt_1p0.gds807
 PIN vccdgt_1p0.gds808
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.418 12.7505 56.458 12.9505 ;
 END
 END vccdgt_1p0.gds808
 PIN vccdgt_1p0.gds809
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.746 12.7505 55.786 12.9505 ;
 END
 END vccdgt_1p0.gds809
 PIN vccdgt_1p0.gds810
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.778 11.011 59.838 11.211 ;
 END
 END vccdgt_1p0.gds810
 PIN vccdgt_1p0.gds811
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.946 11.011 60.006 11.211 ;
 END
 END vccdgt_1p0.gds811
 PIN vccdgt_1p0.gds812
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.106 11.011 59.166 11.211 ;
 END
 END vccdgt_1p0.gds812
 PIN vccdgt_1p0.gds813
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.274 11.011 59.334 11.211 ;
 END
 END vccdgt_1p0.gds813
 PIN vccdgt_1p0.gds814
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.434 11.011 58.494 11.211 ;
 END
 END vccdgt_1p0.gds814
 PIN vccdgt_1p0.gds815
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.602 11.011 58.662 11.211 ;
 END
 END vccdgt_1p0.gds815
 PIN vccdgt_1p0.gds816
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.342 11.011 57.402 11.211 ;
 END
 END vccdgt_1p0.gds816
 PIN vccdgt_1p0.gds817
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.51 11.011 57.57 11.211 ;
 END
 END vccdgt_1p0.gds817
 PIN vccdgt_1p0.gds818
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.67 11.011 56.73 11.211 ;
 END
 END vccdgt_1p0.gds818
 PIN vccdgt_1p0.gds819
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.838 11.011 56.898 11.211 ;
 END
 END vccdgt_1p0.gds819
 PIN vccdgt_1p0.gds820
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.998 11.011 56.058 11.211 ;
 END
 END vccdgt_1p0.gds820
 PIN vccdgt_1p0.gds821
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.166 11.011 56.226 11.211 ;
 END
 END vccdgt_1p0.gds821
 PIN vccdgt_1p0.gds822
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.326 11.011 55.386 11.211 ;
 END
 END vccdgt_1p0.gds822
 PIN vccdgt_1p0.gds823
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.494 11.011 55.554 11.211 ;
 END
 END vccdgt_1p0.gds823
 PIN vccdgt_1p0.gds824
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.922 15.406 59.962 15.606 ;
 END
 END vccdgt_1p0.gds824
 PIN vccdgt_1p0.gds825
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.25 15.406 59.29 15.606 ;
 END
 END vccdgt_1p0.gds825
 PIN vccdgt_1p0.gds826
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.814 15.406 56.854 15.606 ;
 END
 END vccdgt_1p0.gds826
 PIN vccdgt_1p0.gds827
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.142 15.406 56.182 15.606 ;
 END
 END vccdgt_1p0.gds827
 PIN vccdgt_1p0.gds828
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.47 15.406 55.51 15.606 ;
 END
 END vccdgt_1p0.gds828
 PIN vccdgt_1p0.gds829
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.05 13.483 60.09 13.683 ;
 END
 END vccdgt_1p0.gds829
 PIN vccdgt_1p0.gds830
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.73 12.617 59.77 12.817 ;
 END
 END vccdgt_1p0.gds830
 PIN vccdgt_1p0.gds831
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.378 13.483 59.418 13.683 ;
 END
 END vccdgt_1p0.gds831
 PIN vccdgt_1p0.gds832
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.922 11.9905 59.962 12.1905 ;
 END
 END vccdgt_1p0.gds832
 PIN vccdgt_1p0.gds833
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.058 12.617 59.098 12.817 ;
 END
 END vccdgt_1p0.gds833
 PIN vccdgt_1p0.gds834
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.706 13.483 58.746 13.683 ;
 END
 END vccdgt_1p0.gds834
 PIN vccdgt_1p0.gds835
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.25 11.9905 59.29 12.1905 ;
 END
 END vccdgt_1p0.gds835
 PIN vccdgt_1p0.gds836
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.386 12.617 58.426 12.817 ;
 END
 END vccdgt_1p0.gds836
 PIN vccdgt_1p0.gds837
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.034 13.4245 58.074 13.6245 ;
 END
 END vccdgt_1p0.gds837
 PIN vccdgt_1p0.gds838
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.578 11.9905 58.618 12.1905 ;
 END
 END vccdgt_1p0.gds838
 PIN vccdgt_1p0.gds839
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.294 12.617 57.334 12.817 ;
 END
 END vccdgt_1p0.gds839
 PIN vccdgt_1p0.gds840
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.942 13.483 56.982 13.683 ;
 END
 END vccdgt_1p0.gds840
 PIN vccdgt_1p0.gds841
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.486 11.9905 57.526 12.1905 ;
 END
 END vccdgt_1p0.gds841
 PIN vccdgt_1p0.gds842
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.622 12.617 56.662 12.817 ;
 END
 END vccdgt_1p0.gds842
 PIN vccdgt_1p0.gds843
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.27 13.483 56.31 13.683 ;
 END
 END vccdgt_1p0.gds843
 PIN vccdgt_1p0.gds844
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.814 11.9905 56.854 12.1905 ;
 END
 END vccdgt_1p0.gds844
 PIN vccdgt_1p0.gds845
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.95 12.617 55.99 12.817 ;
 END
 END vccdgt_1p0.gds845
 PIN vccdgt_1p0.gds846
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.598 13.483 55.638 13.683 ;
 END
 END vccdgt_1p0.gds846
 PIN vccdgt_1p0.gds847
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.142 11.9905 56.182 12.1905 ;
 END
 END vccdgt_1p0.gds847
 PIN vccdgt_1p0.gds848
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.47 11.9905 55.51 12.1905 ;
 END
 END vccdgt_1p0.gds848
 PIN vccdgt_1p0.gds849
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.578 15.406 58.618 15.606 ;
 END
 END vccdgt_1p0.gds849
 PIN vccdgt_1p0.gds850
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.486 15.406 57.526 15.606 ;
 END
 END vccdgt_1p0.gds850
 PIN vccdgt_1p0.gds851
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.762 13.0135 57.802 13.2135 ;
 END
 END vccdgt_1p0.gds851
 PIN vccdgt_1p0.gds852
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 60.116 15.23 60.172 15.43 ;
 RECT 59.444 15.23 59.5 15.43 ;
 RECT 58.1 15.23 58.156 15.43 ;
 RECT 58.772 15.23 58.828 15.43 ;
 RECT 57.68 15.23 57.736 15.43 ;
 RECT 57.008 15.23 57.064 15.43 ;
 RECT 56.336 15.23 56.392 15.43 ;
 RECT 55.664 15.23 55.72 15.43 ;
 RECT 59.78 12.165 59.836 12.365 ;
 RECT 59.612 12.165 59.668 12.365 ;
 RECT 59.948 12.165 60.004 12.365 ;
 RECT 60.116 12.1635 60.172 12.3635 ;
 RECT 59.108 12.165 59.164 12.365 ;
 RECT 58.94 12.165 58.996 12.365 ;
 RECT 59.276 12.165 59.332 12.365 ;
 RECT 59.444 12.1635 59.5 12.3635 ;
 RECT 58.436 12.165 58.492 12.365 ;
 RECT 58.268 12.165 58.324 12.365 ;
 RECT 58.604 12.165 58.66 12.365 ;
 RECT 58.772 12.1635 58.828 12.3635 ;
 RECT 57.344 12.165 57.4 12.365 ;
 RECT 57.176 12.165 57.232 12.365 ;
 RECT 57.512 12.165 57.568 12.365 ;
 RECT 57.68 12.1635 57.736 12.3635 ;
 RECT 56.672 12.165 56.728 12.365 ;
 RECT 56.504 12.165 56.56 12.365 ;
 RECT 56.84 12.165 56.896 12.365 ;
 RECT 57.008 12.1635 57.064 12.3635 ;
 RECT 56 12.165 56.056 12.365 ;
 RECT 55.832 12.165 55.888 12.365 ;
 RECT 56.168 12.165 56.224 12.365 ;
 RECT 56.336 12.1635 56.392 12.3635 ;
 RECT 55.328 12.165 55.384 12.365 ;
 RECT 55.496 12.165 55.552 12.365 ;
 RECT 55.664 12.1635 55.72 12.3635 ;
 RECT 57.932 13.659 57.988 13.859 ;
 RECT 58.016 13.095 58.072 13.295 ;
 RECT 57.764 13.2495 57.82 13.4495 ;
 RECT 59.78 13.197 59.836 13.397 ;
 RECT 59.612 13.197 59.668 13.397 ;
 RECT 60.116 13.214 60.172 13.414 ;
 RECT 59.948 13.197 60.004 13.397 ;
 RECT 59.108 13.197 59.164 13.397 ;
 RECT 58.94 13.197 58.996 13.397 ;
 RECT 59.444 13.214 59.5 13.414 ;
 RECT 59.276 13.197 59.332 13.397 ;
 RECT 58.436 13.197 58.492 13.397 ;
 RECT 58.268 13.197 58.324 13.397 ;
 RECT 58.1 13.214 58.156 13.414 ;
 RECT 58.772 13.214 58.828 13.414 ;
 RECT 58.604 13.197 58.66 13.397 ;
 RECT 57.344 13.197 57.4 13.397 ;
 RECT 57.176 13.197 57.232 13.397 ;
 RECT 57.68 13.214 57.736 13.414 ;
 RECT 57.512 13.197 57.568 13.397 ;
 RECT 56.672 13.197 56.728 13.397 ;
 RECT 56.504 13.197 56.56 13.397 ;
 RECT 57.008 13.214 57.064 13.414 ;
 RECT 56.84 13.197 56.896 13.397 ;
 RECT 56 13.197 56.056 13.397 ;
 RECT 55.832 13.197 55.888 13.397 ;
 RECT 56.336 13.214 56.392 13.414 ;
 RECT 56.168 13.197 56.224 13.397 ;
 RECT 55.328 13.197 55.384 13.397 ;
 RECT 55.664 13.214 55.72 13.414 ;
 RECT 55.496 13.197 55.552 13.397 ;
 END
 END vccdgt_1p0.gds852
 PIN vccdgt_1p0.gds853
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.97 11.011 63.03 11.211 ;
 END
 END vccdgt_1p0.gds853
 PIN vccdgt_1p0.gds854
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.298 11.011 62.358 11.211 ;
 END
 END vccdgt_1p0.gds854
 PIN vccdgt_1p0.gds855
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.626 11.011 61.686 11.211 ;
 END
 END vccdgt_1p0.gds855
 PIN vccdgt_1p0.gds856
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.954 11.011 61.014 11.211 ;
 END
 END vccdgt_1p0.gds856
 PIN vccdgt_1p0.gds857
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.282 11.011 60.342 11.211 ;
 END
 END vccdgt_1p0.gds857
 PIN vccdgt_1p0.gds858
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.41 13.309 63.45 13.509 ;
 END
 END vccdgt_1p0.gds858
 PIN vccdgt_1p0.gds859
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.886 12.7505 62.926 12.9505 ;
 END
 END vccdgt_1p0.gds859
 PIN vccdgt_1p0.gds860
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.214 12.7505 62.254 12.9505 ;
 END
 END vccdgt_1p0.gds860
 PIN vccdgt_1p0.gds861
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.542 12.7505 61.582 12.9505 ;
 END
 END vccdgt_1p0.gds861
 PIN vccdgt_1p0.gds862
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.87 12.7505 60.91 12.9505 ;
 END
 END vccdgt_1p0.gds862
 PIN vccdgt_1p0.gds863
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.138 11.011 63.198 11.211 ;
 END
 END vccdgt_1p0.gds863
 PIN vccdgt_1p0.gds864
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.306 11.011 63.366 11.211 ;
 END
 END vccdgt_1p0.gds864
 PIN vccdgt_1p0.gds865
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.466 11.011 62.526 11.211 ;
 END
 END vccdgt_1p0.gds865
 PIN vccdgt_1p0.gds866
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.634 11.011 62.694 11.211 ;
 END
 END vccdgt_1p0.gds866
 PIN vccdgt_1p0.gds867
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.794 11.011 61.854 11.211 ;
 END
 END vccdgt_1p0.gds867
 PIN vccdgt_1p0.gds868
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.962 11.011 62.022 11.211 ;
 END
 END vccdgt_1p0.gds868
 PIN vccdgt_1p0.gds869
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.122 11.011 61.182 11.211 ;
 END
 END vccdgt_1p0.gds869
 PIN vccdgt_1p0.gds870
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.29 11.011 61.35 11.211 ;
 END
 END vccdgt_1p0.gds870
 PIN vccdgt_1p0.gds871
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.45 11.011 60.51 11.211 ;
 END
 END vccdgt_1p0.gds871
 PIN vccdgt_1p0.gds872
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.618 11.011 60.678 11.211 ;
 END
 END vccdgt_1p0.gds872
 PIN vccdgt_1p0.gds873
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.498 10.662 64.554 10.862 ;
 END
 END vccdgt_1p0.gds873
 PIN vccdgt_1p0.gds874
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.578 15.003 64.634 15.203 ;
 END
 END vccdgt_1p0.gds874
 PIN vccdgt_1p0.gds875
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.61 15.406 62.65 15.606 ;
 END
 END vccdgt_1p0.gds875
 PIN vccdgt_1p0.gds876
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.938 15.406 61.978 15.606 ;
 END
 END vccdgt_1p0.gds876
 PIN vccdgt_1p0.gds877
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.266 15.406 61.306 15.606 ;
 END
 END vccdgt_1p0.gds877
 PIN vccdgt_1p0.gds878
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.594 15.406 60.634 15.606 ;
 END
 END vccdgt_1p0.gds878
 PIN vccdgt_1p0.gds879
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.09 12.617 63.13 12.817 ;
 END
 END vccdgt_1p0.gds879
 PIN vccdgt_1p0.gds880
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.738 13.483 62.778 13.683 ;
 END
 END vccdgt_1p0.gds880
 PIN vccdgt_1p0.gds881
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.282 11.9905 63.322 12.1905 ;
 END
 END vccdgt_1p0.gds881
 PIN vccdgt_1p0.gds882
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.418 12.617 62.458 12.817 ;
 END
 END vccdgt_1p0.gds882
 PIN vccdgt_1p0.gds883
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.066 13.483 62.106 13.683 ;
 END
 END vccdgt_1p0.gds883
 PIN vccdgt_1p0.gds884
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.61 11.9905 62.65 12.1905 ;
 END
 END vccdgt_1p0.gds884
 PIN vccdgt_1p0.gds885
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.746 12.617 61.786 12.817 ;
 END
 END vccdgt_1p0.gds885
 PIN vccdgt_1p0.gds886
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.394 13.483 61.434 13.683 ;
 END
 END vccdgt_1p0.gds886
 PIN vccdgt_1p0.gds887
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.938 11.9905 61.978 12.1905 ;
 END
 END vccdgt_1p0.gds887
 PIN vccdgt_1p0.gds888
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.074 12.617 61.114 12.817 ;
 END
 END vccdgt_1p0.gds888
 PIN vccdgt_1p0.gds889
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.722 13.483 60.762 13.683 ;
 END
 END vccdgt_1p0.gds889
 PIN vccdgt_1p0.gds890
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.266 11.9905 61.306 12.1905 ;
 END
 END vccdgt_1p0.gds890
 PIN vccdgt_1p0.gds891
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.402 12.617 60.442 12.817 ;
 END
 END vccdgt_1p0.gds891
 PIN vccdgt_1p0.gds892
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.594 11.9905 60.634 12.1905 ;
 END
 END vccdgt_1p0.gds892
 PIN vccdgt_1p0.gds893
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.658 10.8945 64.714 11.0945 ;
 END
 END vccdgt_1p0.gds893
 PIN vccdgt_1p0.gds894
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.078 11.224 64.134 11.424 ;
 END
 END vccdgt_1p0.gds894
 PIN vccdgt_1p0.gds895
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.078 14.7305 64.134 14.9305 ;
 END
 END vccdgt_1p0.gds895
 PIN vccdgt_1p0.gds896
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.318 13.189 64.394 13.389 ;
 END
 END vccdgt_1p0.gds896
 PIN vccdgt_1p0.gds897
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.158 13.803 65.234 14.003 ;
 END
 END vccdgt_1p0.gds897
 PIN vccdgt_1p0.gds898
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.282 15.406 63.322 15.606 ;
 END
 END vccdgt_1p0.gds898
 PIN vccdgt_1p0.gds899
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.834 10.478 63.874 10.678 ;
 END
 END vccdgt_1p0.gds899
 PIN vccdgt_1p0.gds900
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.558 13.446 63.618 13.646 ;
 END
 END vccdgt_1p0.gds900
 PIN vccdgt_1p0.gds901
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 63.896 15.091 63.952 15.291 ;
 RECT 64.232 15.127 64.288 15.309 ;
 RECT 64.568 15.127 64.624 15.309 ;
 RECT 64.904 15.127 64.96 15.309 ;
 RECT 63.896 15.37 63.952 15.57 ;
 RECT 64.736 15.37 64.792 15.57 ;
 RECT 64.4 15.3035 64.456 15.5035 ;
 RECT 64.064 15.4105 64.12 15.6105 ;
 RECT 65.072 15.2705 65.128 15.4705 ;
 RECT 63.476 15.23 63.532 15.43 ;
 RECT 62.804 15.23 62.86 15.43 ;
 RECT 62.132 15.23 62.188 15.43 ;
 RECT 61.46 15.23 61.516 15.43 ;
 RECT 60.788 15.23 60.844 15.43 ;
 RECT 64.568 14.007 64.624 14.189 ;
 RECT 64.4 13.989 64.456 14.189 ;
 RECT 64.904 14.007 64.96 14.189 ;
 RECT 64.652 12.682 64.708 12.882 ;
 RECT 64.232 12.682 64.288 12.882 ;
 RECT 63.812 12.403 63.868 12.603 ;
 RECT 64.568 12.439 64.624 12.621 ;
 RECT 64.4 12.439 64.456 12.621 ;
 RECT 64.232 12.439 64.288 12.621 ;
 RECT 65.072 12.542 65.128 12.742 ;
 RECT 64.904 12.439 64.96 12.621 ;
 RECT 63.812 11.337 63.868 11.537 ;
 RECT 64.232 11.319 64.288 11.501 ;
 RECT 64.568 11.319 64.624 11.501 ;
 RECT 64.4 11.319 64.456 11.501 ;
 RECT 65.072 11.319 65.128 11.501 ;
 RECT 64.904 11.319 64.96 11.501 ;
 RECT 64.064 11.058 64.12 11.258 ;
 RECT 65.072 11.058 65.128 11.258 ;
 RECT 64.736 11.058 64.792 11.258 ;
 RECT 64.4 11.058 64.456 11.258 ;
 RECT 63.812 11.059 63.868 11.259 ;
 RECT 64.652 13.676 64.708 13.876 ;
 RECT 64.232 13.886 64.288 14.086 ;
 RECT 65.072 13.7925 65.128 13.9925 ;
 RECT 64.064 13.634 64.12 13.834 ;
 RECT 63.728 14.1515 63.784 14.3515 ;
 RECT 63.14 12.165 63.196 12.365 ;
 RECT 62.972 12.165 63.028 12.365 ;
 RECT 63.308 12.165 63.364 12.365 ;
 RECT 63.476 12.1635 63.532 12.3635 ;
 RECT 62.468 12.165 62.524 12.365 ;
 RECT 62.3 12.165 62.356 12.365 ;
 RECT 62.636 12.165 62.692 12.365 ;
 RECT 62.804 12.1635 62.86 12.3635 ;
 RECT 61.796 12.165 61.852 12.365 ;
 RECT 61.628 12.165 61.684 12.365 ;
 RECT 61.964 12.165 62.02 12.365 ;
 RECT 62.132 12.1635 62.188 12.3635 ;
 RECT 61.124 12.165 61.18 12.365 ;
 RECT 60.956 12.165 61.012 12.365 ;
 RECT 61.292 12.165 61.348 12.365 ;
 RECT 61.46 12.1635 61.516 12.3635 ;
 RECT 60.452 12.165 60.508 12.365 ;
 RECT 60.62 12.165 60.676 12.365 ;
 RECT 60.788 12.1635 60.844 12.3635 ;
 RECT 60.284 12.165 60.34 12.365 ;
 RECT 63.14 13.197 63.196 13.397 ;
 RECT 62.972 13.197 63.028 13.397 ;
 RECT 63.476 13.214 63.532 13.414 ;
 RECT 63.308 13.197 63.364 13.397 ;
 RECT 62.468 13.197 62.524 13.397 ;
 RECT 62.3 13.197 62.356 13.397 ;
 RECT 62.804 13.214 62.86 13.414 ;
 RECT 62.636 13.197 62.692 13.397 ;
 RECT 61.796 13.197 61.852 13.397 ;
 RECT 61.628 13.197 61.684 13.397 ;
 RECT 62.132 13.214 62.188 13.414 ;
 RECT 61.964 13.197 62.02 13.397 ;
 RECT 61.124 13.197 61.18 13.397 ;
 RECT 60.956 13.197 61.012 13.397 ;
 RECT 61.46 13.214 61.516 13.414 ;
 RECT 61.292 13.197 61.348 13.397 ;
 RECT 60.452 13.197 60.508 13.397 ;
 RECT 60.788 13.214 60.844 13.414 ;
 RECT 60.62 13.197 60.676 13.397 ;
 RECT 60.284 13.197 60.34 13.397 ;
 END
 END vccdgt_1p0.gds901
 PIN vccdgt_1p0.gds902
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.194 11.011 70.254 11.211 ;
 END
 END vccdgt_1p0.gds902
 PIN vccdgt_1p0.gds903
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.522 11.011 69.582 11.211 ;
 END
 END vccdgt_1p0.gds903
 PIN vccdgt_1p0.gds904
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.69 11.011 69.75 11.211 ;
 END
 END vccdgt_1p0.gds904
 PIN vccdgt_1p0.gds905
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.858 11.011 69.918 11.211 ;
 END
 END vccdgt_1p0.gds905
 PIN vccdgt_1p0.gds906
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.11 12.7505 70.15 12.9505 ;
 END
 END vccdgt_1p0.gds906
 PIN vccdgt_1p0.gds907
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.438 12.7505 69.478 12.9505 ;
 END
 END vccdgt_1p0.gds907
 PIN vccdgt_1p0.gds908
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.174 13.1425 68.23 13.3425 ;
 END
 END vccdgt_1p0.gds908
 PIN vccdgt_1p0.gds909
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.994 12.5175 68.05 12.7175 ;
 END
 END vccdgt_1p0.gds909
 PIN vccdgt_1p0.gds910
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 10.502 67.726 10.702 ;
 END
 END vccdgt_1p0.gds910
 PIN vccdgt_1p0.gds911
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.022 14.062 67.082 14.262 ;
 END
 END vccdgt_1p0.gds911
 PIN vccdgt_1p0.gds912
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.49 13.268 67.546 13.468 ;
 END
 END vccdgt_1p0.gds912
 PIN vccdgt_1p0.gds913
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.642 12.617 69.682 12.817 ;
 END
 END vccdgt_1p0.gds913
 PIN vccdgt_1p0.gds914
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 13.374 68.89 13.574 ;
 END
 END vccdgt_1p0.gds914
 PIN vccdgt_1p0.gds915
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.342 12.527 66.382 12.727 ;
 END
 END vccdgt_1p0.gds915
 PIN vccdgt_1p0.gds916
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.922 11.95 65.962 12.15 ;
 END
 END vccdgt_1p0.gds916
 PIN vccdgt_1p0.gds917
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.338 12.7505 65.394 12.9505 ;
 END
 END vccdgt_1p0.gds917
 PIN vccdgt_1p0.gds918
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.014 11.6505 69.054 11.8505 ;
 END
 END vccdgt_1p0.gds918
 PIN vccdgt_1p0.gds919
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.678 12.3155 66.738 12.5155 ;
 END
 END vccdgt_1p0.gds919
 PIN vccdgt_1p0.gds920
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.754 11.025 68.81 11.225 ;
 END
 END vccdgt_1p0.gds920
 PIN vccdgt_1p0.gds921
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.962 13.483 70.002 13.683 ;
 END
 END vccdgt_1p0.gds921
 PIN vccdgt_1p0.gds922
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.834 11.9905 69.874 12.1905 ;
 END
 END vccdgt_1p0.gds922
 PIN vccdgt_1p0.gds923
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.494 13.2505 68.57 13.4505 ;
 END
 END vccdgt_1p0.gds923
 PIN vccdgt_1p0.gds924
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.83 12.968 67.89 13.168 ;
 END
 END vccdgt_1p0.gds924
 PIN vccdgt_1p0.gds925
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.47 14.213 66.51 14.413 ;
 END
 END vccdgt_1p0.gds925
 PIN vccdgt_1p0.gds926
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.758 13.638 65.814 13.838 ;
 END
 END vccdgt_1p0.gds926
 PIN vccdgt_1p0.gds927
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.27 13.2825 69.33 13.4825 ;
 END
 END vccdgt_1p0.gds927
 PIN vccdgt_1p0.gds928
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.334 13.0715 68.39 13.2715 ;
 END
 END vccdgt_1p0.gds928
 PIN vccdgt_1p0.gds929
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.114 14.05 66.154 14.25 ;
 END
 END vccdgt_1p0.gds929
 PIN vccdgt_1p0.gds930
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.186 14.161 67.232 14.361 ;
 END
 END vccdgt_1p0.gds930
 PIN vccdgt_1p0.gds931
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.834 15.406 69.874 15.606 ;
 END
 END vccdgt_1p0.gds931
 PIN vccdgt_1p0.gds932
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 65.24 15.127 65.296 15.309 ;
 RECT 66.248 15.09 66.304 15.29 ;
 RECT 65.912 15.09 65.968 15.29 ;
 RECT 66.584 15.09 66.64 15.29 ;
 RECT 67.844 15.109 67.9 15.309 ;
 RECT 67.424 15.127 67.48 15.309 ;
 RECT 68.936 15.091 68.992 15.291 ;
 RECT 66.416 15.37 66.472 15.57 ;
 RECT 66.08 15.37 66.136 15.57 ;
 RECT 67.088 15.37 67.144 15.57 ;
 RECT 66.752 15.37 66.808 15.57 ;
 RECT 67.424 15.37 67.48 15.57 ;
 RECT 68.684 15.23 68.74 15.43 ;
 RECT 68.348 15.351 68.404 15.533 ;
 RECT 68.936 15.369 68.992 15.569 ;
 RECT 69.356 15.23 69.412 15.43 ;
 RECT 70.028 15.23 70.084 15.43 ;
 RECT 65.408 14.007 65.464 14.189 ;
 RECT 65.24 14.007 65.296 14.189 ;
 RECT 66.248 14.026 66.304 14.226 ;
 RECT 65.912 14.026 65.968 14.226 ;
 RECT 65.744 14.007 65.8 14.189 ;
 RECT 66.584 14.026 66.64 14.226 ;
 RECT 67.088 14.007 67.144 14.189 ;
 RECT 66.92 14.007 66.976 14.189 ;
 RECT 67.844 14.007 67.9 14.189 ;
 RECT 67.676 14.007 67.732 14.189 ;
 RECT 67.508 14.007 67.564 14.189 ;
 RECT 68.516 14.007 68.572 14.189 ;
 RECT 68.348 14.007 68.404 14.189 ;
 RECT 69.272 14.064 69.328 14.264 ;
 RECT 66.332 12.682 66.388 12.882 ;
 RECT 65.996 12.682 66.052 12.882 ;
 RECT 67.256 12.679 67.312 12.843 ;
 RECT 66.668 12.682 66.724 12.882 ;
 RECT 67.004 12.672 67.06 12.843 ;
 RECT 68.684 12.681 68.74 12.881 ;
 RECT 65.492 12.542 65.548 12.742 ;
 RECT 65.24 12.439 65.296 12.621 ;
 RECT 65.996 12.402 66.052 12.602 ;
 RECT 65.828 12.542 65.884 12.742 ;
 RECT 67.088 12.439 67.144 12.621 ;
 RECT 66.92 12.439 66.976 12.621 ;
 RECT 66.752 12.439 66.808 12.621 ;
 RECT 66.584 12.439 66.64 12.621 ;
 RECT 67.76 12.403 67.816 12.603 ;
 RECT 67.34 12.441 67.396 12.621 ;
 RECT 68.684 12.403 68.74 12.603 ;
 RECT 68.432 12.3615 68.488 12.5615 ;
 RECT 68.264 12.3615 68.32 12.5615 ;
 RECT 68.096 12.402 68.152 12.602 ;
 RECT 68.936 12.403 68.992 12.603 ;
 RECT 65.492 11.319 65.548 11.501 ;
 RECT 65.24 11.319 65.296 11.501 ;
 RECT 65.996 11.319 66.052 11.501 ;
 RECT 65.828 11.301 65.884 11.501 ;
 RECT 66.92 11.301 66.976 11.501 ;
 RECT 66.752 11.301 66.808 11.501 ;
 RECT 66.584 11.301 66.64 11.501 ;
 RECT 67.844 11.338 67.9 11.538 ;
 RECT 67.676 11.301 67.732 11.501 ;
 RECT 67.508 11.301 67.564 11.501 ;
 RECT 68.684 11.301 68.74 11.501 ;
 RECT 69.02 11.337 69.076 11.537 ;
 RECT 66.08 11.058 66.136 11.258 ;
 RECT 65.744 11.058 65.8 11.258 ;
 RECT 67.76 11.058 67.816 11.258 ;
 RECT 68.096 11.058 68.152 11.258 ;
 RECT 66.332 13.746 66.388 13.946 ;
 RECT 65.996 13.746 66.052 13.946 ;
 RECT 65.828 13.783 65.884 13.965 ;
 RECT 67.256 13.8845 67.312 14.0845 ;
 RECT 66.668 13.746 66.724 13.946 ;
 RECT 67.004 13.785 67.06 13.951 ;
 RECT 65.408 15.249 65.464 15.449 ;
 RECT 65.408 10.988 65.464 11.188 ;
 RECT 70.196 12.165 70.252 12.365 ;
 RECT 69.692 12.165 69.748 12.365 ;
 RECT 69.524 12.165 69.58 12.365 ;
 RECT 69.86 12.165 69.916 12.365 ;
 RECT 70.028 12.1635 70.084 12.3635 ;
 RECT 68.18 12.752 68.236 12.952 ;
 RECT 67.676 12.752 67.732 12.952 ;
 RECT 68.852 11.267 68.908 11.467 ;
 RECT 68.096 11.408 68.152 11.608 ;
 RECT 68.432 11.291 68.488 11.491 ;
 RECT 68.264 11.408 68.32 11.608 ;
 RECT 67.424 10.988 67.48 11.188 ;
 RECT 67.088 11.1275 67.144 11.3275 ;
 RECT 67.34 11.2685 67.396 11.4685 ;
 RECT 67.004 15.02 67.06 15.22 ;
 RECT 68.432 15.02 68.488 15.22 ;
 RECT 68.264 15.02 68.32 15.22 ;
 RECT 67.172 15.09 67.228 15.29 ;
 RECT 65.66 15.2025 65.716 15.4025 ;
 RECT 67.676 15.127 67.732 15.309 ;
 RECT 68.6 15.239 68.656 15.439 ;
 RECT 68.096 15.351 68.152 15.533 ;
 RECT 69.188 14.5165 69.244 14.7165 ;
 RECT 67.76 13.676 67.816 13.876 ;
 RECT 68.684 13.7265 68.74 13.9265 ;
 RECT 68.264 13.676 68.32 13.876 ;
 RECT 65.492 13.676 65.548 13.876 ;
 RECT 70.196 13.197 70.252 13.397 ;
 RECT 69.692 13.197 69.748 13.397 ;
 RECT 69.524 13.197 69.58 13.397 ;
 RECT 69.356 13.214 69.412 13.414 ;
 RECT 70.028 13.214 70.084 13.414 ;
 RECT 69.86 13.197 69.916 13.397 ;
 END
 END vccdgt_1p0.gds932
 PIN vccdgt_1p0.gds933
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.226 11.011 74.286 11.211 ;
 END
 END vccdgt_1p0.gds933
 PIN vccdgt_1p0.gds934
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.554 11.011 73.614 11.211 ;
 END
 END vccdgt_1p0.gds934
 PIN vccdgt_1p0.gds935
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.882 11.011 72.942 11.211 ;
 END
 END vccdgt_1p0.gds935
 PIN vccdgt_1p0.gds936
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.21 11.011 72.27 11.211 ;
 END
 END vccdgt_1p0.gds936
 PIN vccdgt_1p0.gds937
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.538 11.011 71.598 11.211 ;
 END
 END vccdgt_1p0.gds937
 PIN vccdgt_1p0.gds938
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.866 11.011 70.926 11.211 ;
 END
 END vccdgt_1p0.gds938
 PIN vccdgt_1p0.gds939
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.394 11.011 74.454 11.211 ;
 END
 END vccdgt_1p0.gds939
 PIN vccdgt_1p0.gds940
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.562 11.011 74.622 11.211 ;
 END
 END vccdgt_1p0.gds940
 PIN vccdgt_1p0.gds941
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.722 11.011 73.782 11.211 ;
 END
 END vccdgt_1p0.gds941
 PIN vccdgt_1p0.gds942
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.89 11.011 73.95 11.211 ;
 END
 END vccdgt_1p0.gds942
 PIN vccdgt_1p0.gds943
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.05 11.011 73.11 11.211 ;
 END
 END vccdgt_1p0.gds943
 PIN vccdgt_1p0.gds944
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.218 11.011 73.278 11.211 ;
 END
 END vccdgt_1p0.gds944
 PIN vccdgt_1p0.gds945
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.378 11.011 72.438 11.211 ;
 END
 END vccdgt_1p0.gds945
 PIN vccdgt_1p0.gds946
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.546 11.011 72.606 11.211 ;
 END
 END vccdgt_1p0.gds946
 PIN vccdgt_1p0.gds947
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.706 11.011 71.766 11.211 ;
 END
 END vccdgt_1p0.gds947
 PIN vccdgt_1p0.gds948
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.874 11.011 71.934 11.211 ;
 END
 END vccdgt_1p0.gds948
 PIN vccdgt_1p0.gds949
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.034 11.011 71.094 11.211 ;
 END
 END vccdgt_1p0.gds949
 PIN vccdgt_1p0.gds950
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.202 11.011 71.262 11.211 ;
 END
 END vccdgt_1p0.gds950
 PIN vccdgt_1p0.gds951
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.362 11.011 70.422 11.211 ;
 END
 END vccdgt_1p0.gds951
 PIN vccdgt_1p0.gds952
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.53 11.011 70.59 11.211 ;
 END
 END vccdgt_1p0.gds952
 PIN vccdgt_1p0.gds953
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.666 13.309 74.706 13.509 ;
 END
 END vccdgt_1p0.gds953
 PIN vccdgt_1p0.gds954
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.142 12.7505 74.182 12.9505 ;
 END
 END vccdgt_1p0.gds954
 PIN vccdgt_1p0.gds955
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.47 12.7505 73.51 12.9505 ;
 END
 END vccdgt_1p0.gds955
 PIN vccdgt_1p0.gds956
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.798 12.7505 72.838 12.9505 ;
 END
 END vccdgt_1p0.gds956
 PIN vccdgt_1p0.gds957
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.126 12.7505 72.166 12.9505 ;
 END
 END vccdgt_1p0.gds957
 PIN vccdgt_1p0.gds958
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.454 12.7505 71.494 12.9505 ;
 END
 END vccdgt_1p0.gds958
 PIN vccdgt_1p0.gds959
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.782 12.7505 70.822 12.9505 ;
 END
 END vccdgt_1p0.gds959
 PIN vccdgt_1p0.gds960
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.538 15.406 74.578 15.606 ;
 END
 END vccdgt_1p0.gds960
 PIN vccdgt_1p0.gds961
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.866 15.406 73.906 15.606 ;
 END
 END vccdgt_1p0.gds961
 PIN vccdgt_1p0.gds962
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.194 15.406 73.234 15.606 ;
 END
 END vccdgt_1p0.gds962
 PIN vccdgt_1p0.gds963
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.522 15.406 72.562 15.606 ;
 END
 END vccdgt_1p0.gds963
 PIN vccdgt_1p0.gds964
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.85 15.406 71.89 15.606 ;
 END
 END vccdgt_1p0.gds964
 PIN vccdgt_1p0.gds965
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.178 15.406 71.218 15.606 ;
 END
 END vccdgt_1p0.gds965
 PIN vccdgt_1p0.gds966
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.506 15.406 70.546 15.606 ;
 END
 END vccdgt_1p0.gds966
 PIN vccdgt_1p0.gds967
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.346 12.617 74.386 12.817 ;
 END
 END vccdgt_1p0.gds967
 PIN vccdgt_1p0.gds968
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.994 13.483 74.034 13.683 ;
 END
 END vccdgt_1p0.gds968
 PIN vccdgt_1p0.gds969
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.538 11.9905 74.578 12.1905 ;
 END
 END vccdgt_1p0.gds969
 PIN vccdgt_1p0.gds970
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.674 12.617 73.714 12.817 ;
 END
 END vccdgt_1p0.gds970
 PIN vccdgt_1p0.gds971
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.322 13.483 73.362 13.683 ;
 END
 END vccdgt_1p0.gds971
 PIN vccdgt_1p0.gds972
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.866 11.9905 73.906 12.1905 ;
 END
 END vccdgt_1p0.gds972
 PIN vccdgt_1p0.gds973
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.002 12.617 73.042 12.817 ;
 END
 END vccdgt_1p0.gds973
 PIN vccdgt_1p0.gds974
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.65 13.483 72.69 13.683 ;
 END
 END vccdgt_1p0.gds974
 PIN vccdgt_1p0.gds975
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.194 11.9905 73.234 12.1905 ;
 END
 END vccdgt_1p0.gds975
 PIN vccdgt_1p0.gds976
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.33 12.617 72.37 12.817 ;
 END
 END vccdgt_1p0.gds976
 PIN vccdgt_1p0.gds977
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.978 13.483 72.018 13.683 ;
 END
 END vccdgt_1p0.gds977
 PIN vccdgt_1p0.gds978
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.522 11.9905 72.562 12.1905 ;
 END
 END vccdgt_1p0.gds978
 PIN vccdgt_1p0.gds979
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.658 12.617 71.698 12.817 ;
 END
 END vccdgt_1p0.gds979
 PIN vccdgt_1p0.gds980
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.306 13.483 71.346 13.683 ;
 END
 END vccdgt_1p0.gds980
 PIN vccdgt_1p0.gds981
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.85 11.9905 71.89 12.1905 ;
 END
 END vccdgt_1p0.gds981
 PIN vccdgt_1p0.gds982
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.986 12.617 71.026 12.817 ;
 END
 END vccdgt_1p0.gds982
 PIN vccdgt_1p0.gds983
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.634 13.483 70.674 13.683 ;
 END
 END vccdgt_1p0.gds983
 PIN vccdgt_1p0.gds984
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.178 11.9905 71.218 12.1905 ;
 END
 END vccdgt_1p0.gds984
 PIN vccdgt_1p0.gds985
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.314 12.617 70.354 12.817 ;
 END
 END vccdgt_1p0.gds985
 PIN vccdgt_1p0.gds986
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.506 11.9905 70.546 12.1905 ;
 END
 END vccdgt_1p0.gds986
 PIN vccdgt_1p0.gds987
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 74.732 15.23 74.788 15.43 ;
 RECT 74.06 15.23 74.116 15.43 ;
 RECT 73.388 15.23 73.444 15.43 ;
 RECT 72.716 15.23 72.772 15.43 ;
 RECT 72.044 15.23 72.1 15.43 ;
 RECT 71.372 15.23 71.428 15.43 ;
 RECT 70.7 15.23 70.756 15.43 ;
 RECT 74.396 12.165 74.452 12.365 ;
 RECT 74.228 12.165 74.284 12.365 ;
 RECT 74.564 12.165 74.62 12.365 ;
 RECT 74.732 12.1635 74.788 12.3635 ;
 RECT 73.724 12.165 73.78 12.365 ;
 RECT 73.556 12.165 73.612 12.365 ;
 RECT 73.892 12.165 73.948 12.365 ;
 RECT 74.06 12.1635 74.116 12.3635 ;
 RECT 73.052 12.165 73.108 12.365 ;
 RECT 72.884 12.165 72.94 12.365 ;
 RECT 73.22 12.165 73.276 12.365 ;
 RECT 73.388 12.1635 73.444 12.3635 ;
 RECT 72.38 12.165 72.436 12.365 ;
 RECT 72.212 12.165 72.268 12.365 ;
 RECT 72.548 12.165 72.604 12.365 ;
 RECT 72.716 12.1635 72.772 12.3635 ;
 RECT 71.708 12.165 71.764 12.365 ;
 RECT 71.54 12.165 71.596 12.365 ;
 RECT 71.876 12.165 71.932 12.365 ;
 RECT 72.044 12.1635 72.1 12.3635 ;
 RECT 71.036 12.165 71.092 12.365 ;
 RECT 70.868 12.165 70.924 12.365 ;
 RECT 71.204 12.165 71.26 12.365 ;
 RECT 71.372 12.1635 71.428 12.3635 ;
 RECT 70.364 12.165 70.42 12.365 ;
 RECT 70.532 12.165 70.588 12.365 ;
 RECT 70.7 12.1635 70.756 12.3635 ;
 RECT 74.396 13.197 74.452 13.397 ;
 RECT 74.228 13.197 74.284 13.397 ;
 RECT 74.732 13.214 74.788 13.414 ;
 RECT 74.564 13.197 74.62 13.397 ;
 RECT 73.724 13.197 73.78 13.397 ;
 RECT 73.556 13.197 73.612 13.397 ;
 RECT 74.06 13.214 74.116 13.414 ;
 RECT 73.892 13.197 73.948 13.397 ;
 RECT 73.052 13.197 73.108 13.397 ;
 RECT 72.884 13.197 72.94 13.397 ;
 RECT 73.388 13.214 73.444 13.414 ;
 RECT 73.22 13.197 73.276 13.397 ;
 RECT 72.38 13.197 72.436 13.397 ;
 RECT 72.212 13.197 72.268 13.397 ;
 RECT 72.716 13.214 72.772 13.414 ;
 RECT 72.548 13.197 72.604 13.397 ;
 RECT 71.708 13.197 71.764 13.397 ;
 RECT 71.54 13.197 71.596 13.397 ;
 RECT 72.044 13.214 72.1 13.414 ;
 RECT 71.876 13.197 71.932 13.397 ;
 RECT 71.036 13.197 71.092 13.397 ;
 RECT 70.868 13.197 70.924 13.397 ;
 RECT 71.372 13.214 71.428 13.414 ;
 RECT 71.204 13.197 71.26 13.397 ;
 RECT 70.364 13.197 70.42 13.397 ;
 RECT 70.7 13.214 70.756 13.414 ;
 RECT 70.532 13.197 70.588 13.397 ;
 END
 END vccdgt_1p0.gds987
 PIN vccdgt_1p0.gds988
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 17.344 0.654 17.544 ;
 END
 END vccdgt_1p0.gds988
 PIN vccdgt_1p0.gds989
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 19.343 0.654 19.543 ;
 END
 END vccdgt_1p0.gds989
 PIN vccdgt_1p0.gds990
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.454 17.902 0.494 18.102 ;
 END
 END vccdgt_1p0.gds990
 PIN vccdgt_1p0.gds991
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.566 18.0745 1.622 18.2745 ;
 END
 END vccdgt_1p0.gds991
 PIN vccdgt_1p0.gds992
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.742 18.126 0.788 18.326 ;
 END
 END vccdgt_1p0.gds992
 PIN vccdgt_1p0.gds993
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.114 17.847 1.154 18.047 ;
 END
 END vccdgt_1p0.gds993
 PIN vccdgt_1p0.gds994
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.966 18.064 1.026 18.264 ;
 END
 END vccdgt_1p0.gds994
 PIN vccdgt_1p0.gds995
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.986 18.7015 2.042 18.9015 ;
 END
 END vccdgt_1p0.gds995
 PIN vccdgt_1p0.gds996
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.326 18.175 2.382 18.375 ;
 END
 END vccdgt_1p0.gds996
 PIN vccdgt_1p0.gds997
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.806 18.137 1.882 18.337 ;
 END
 END vccdgt_1p0.gds997
 PIN vccdgt_1p0.gds998
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.166 20.3885 3.206 20.5885 ;
 END
 END vccdgt_1p0.gds998
 PIN vccdgt_1p0.gds999
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.646 17.7935 2.722 17.9935 ;
 END
 END vccdgt_1p0.gds999
 PIN vccdgt_1p0.gds1000
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.098 20.2255 5.138 20.4255 ;
 END
 END vccdgt_1p0.gds1000
 PIN vccdgt_1p0.gds1001
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.634 17.98 4.674 18.18 ;
 END
 END vccdgt_1p0.gds1001
 PIN vccdgt_1p0.gds1002
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.478 17.5525 3.538 17.7525 ;
 END
 END vccdgt_1p0.gds1002
 PIN vccdgt_1p0.gds1003
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.69 16.745 3.73 16.945 ;
 END
 END vccdgt_1p0.gds1003
 PIN vccdgt_1p0.gds1004
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.09 20.088 4.13 20.288 ;
 END
 END vccdgt_1p0.gds1004
 PIN vccdgt_1p0.gds1005
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.906 20.061 4.946 20.261 ;
 END
 END vccdgt_1p0.gds1005
 PIN vccdgt_1p0.gds1006
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.362 17.772 4.418 17.972 ;
 END
 END vccdgt_1p0.gds1006
 PIN vccdgt_1p0.gds1007
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.762 18.154 4.818 18.354 ;
 END
 END vccdgt_1p0.gds1007
 PIN vccdgt_1p0.gds1008
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.486 17.854 2.542 18.054 ;
 END
 END vccdgt_1p0.gds1008
 PIN vccdgt_1p0.gds1009
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 3.248 18.055 3.304 18.219 ;
 RECT 3.752 18.055 3.808 18.219 ;
 RECT 4.004 18.055 4.06 18.219 ;
 RECT 1.988 18.057 2.044 18.257 ;
 RECT 2.492 18.057 2.548 18.257 ;
 RECT 2.24 18.057 2.296 18.257 ;
 RECT 2.996 18.057 3.052 18.257 ;
 RECT 2.744 18.057 2.8 18.257 ;
 RECT 1.568 18.058 1.624 18.258 ;
 RECT 1.4 18.058 1.456 18.258 ;
 RECT 0.896 18.058 0.952 18.258 ;
 RECT 0.56 18.0985 0.616 18.2985 ;
 RECT 4.424 18.057 4.48 18.257 ;
 RECT 4.928 18.039 4.984 18.221 ;
 RECT 3.5 16.471 3.556 16.653 ;
 RECT 0.896 16.434 0.952 16.634 ;
 RECT 0.56 16.434 0.616 16.634 ;
 RECT 1.568 16.434 1.624 16.634 ;
 RECT 1.4 16.434 1.456 16.634 ;
 RECT 2.576 16.434 2.632 16.634 ;
 RECT 2.156 16.434 2.212 16.634 ;
 RECT 1.988 16.434 2.044 16.634 ;
 RECT 4.928 16.471 4.984 16.653 ;
 RECT 3.668 16.5725 3.724 16.7725 ;
 RECT 3.248 16.574 3.304 16.774 ;
 RECT 3.5 16.695 3.556 16.877 ;
 RECT 4.088 16.574 4.144 16.774 ;
 RECT 3.92 16.574 3.976 16.774 ;
 RECT 0.896 16.714 0.952 16.914 ;
 RECT 0.56 16.714 0.616 16.914 ;
 RECT 1.568 16.714 1.624 16.914 ;
 RECT 1.4 16.714 1.456 16.914 ;
 RECT 2.408 16.695 2.464 16.875 ;
 RECT 1.232 19.62 1.288 19.82 ;
 RECT 1.568 19.635 1.624 19.835 ;
 RECT 1.82 19.635 1.876 19.835 ;
 RECT 2.072 19.749 2.128 19.929 ;
 RECT 2.996 19.747 3.052 19.929 ;
 RECT 3.164 19.747 3.22 19.923 ;
 RECT 2.492 19.2485 2.548 19.4485 ;
 RECT 0.812 19.653 0.868 19.853 ;
 RECT 0.644 19.653 0.7 19.853 ;
 RECT 0.98 19.653 1.036 19.853 ;
 RECT 4.088 19.1975 4.144 19.3975 ;
 RECT 4.676 19.1975 4.732 19.3975 ;
 RECT 4.424 19.1975 4.48 19.3975 ;
 RECT 5.012 19.1975 5.068 19.3975 ;
 RECT 4.844 19.1975 4.9 19.3975 ;
 RECT 2.156 16.784 2.212 16.984 ;
 RECT 1.988 16.784 2.044 16.984 ;
 RECT 2.996 16.713 3.052 16.913 ;
 RECT 2.744 16.713 2.8 16.913 ;
 RECT 5.18 16.574 5.236 16.774 ;
 RECT 4.424 16.5725 4.48 16.7725 ;
 RECT 4.928 16.695 4.984 16.877 ;
 RECT 4.676 16.574 4.732 16.774 ;
 RECT 3.668 17.815 3.724 17.997 ;
 RECT 3.248 17.779 3.304 17.979 ;
 RECT 3.5 17.9165 3.556 18.1165 ;
 RECT 4.088 17.778 4.144 17.978 ;
 RECT 3.92 17.778 3.976 17.978 ;
 RECT 0.896 17.778 0.952 17.978 ;
 RECT 0.56 17.778 0.616 17.978 ;
 RECT 1.568 17.778 1.624 17.978 ;
 RECT 1.4 17.778 1.456 17.978 ;
 RECT 2.408 17.778 2.464 17.978 ;
 RECT 2.24 17.778 2.296 17.978 ;
 RECT 2.072 17.778 2.128 17.978 ;
 RECT 2.996 17.779 3.052 17.979 ;
 RECT 2.744 17.779 2.8 17.979 ;
 RECT 4.424 17.779 4.48 17.979 ;
 RECT 4.928 17.815 4.984 17.997 ;
 RECT 4.676 17.918 4.732 18.118 ;
 RECT 5.18 17.918 5.236 18.118 ;
 END
 END vccdgt_1p0.gds1009
 PIN vccdgt_1p0.gds1010
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.714 15.679 9.754 15.879 ;
 END
 END vccdgt_1p0.gds1010
 PIN vccdgt_1p0.gds1011
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.042 15.679 9.082 15.879 ;
 END
 END vccdgt_1p0.gds1011
 PIN vccdgt_1p0.gds1012
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.37 15.679 8.41 15.879 ;
 END
 END vccdgt_1p0.gds1012
 PIN vccdgt_1p0.gds1013
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.698 15.679 7.738 15.879 ;
 END
 END vccdgt_1p0.gds1013
 PIN vccdgt_1p0.gds1014
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.626 18.602 5.666 18.802 ;
 END
 END vccdgt_1p0.gds1014
 PIN vccdgt_1p0.gds1015
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.026 15.679 7.066 15.879 ;
 END
 END vccdgt_1p0.gds1015
 PIN vccdgt_1p0.gds1016
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.33 18.739 6.37 18.939 ;
 END
 END vccdgt_1p0.gds1016
 PIN vccdgt_1p0.gds1017
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.966 17.5555 10.026 17.7555 ;
 END
 END vccdgt_1p0.gds1017
 PIN vccdgt_1p0.gds1018
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.294 17.5555 9.354 17.7555 ;
 END
 END vccdgt_1p0.gds1018
 PIN vccdgt_1p0.gds1019
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.622 17.5555 8.682 17.7555 ;
 END
 END vccdgt_1p0.gds1019
 PIN vccdgt_1p0.gds1020
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.95 17.5555 8.01 17.7555 ;
 END
 END vccdgt_1p0.gds1020
 PIN vccdgt_1p0.gds1021
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.278 17.5555 7.338 17.7555 ;
 END
 END vccdgt_1p0.gds1021
 PIN vccdgt_1p0.gds1022
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.862 18.081 6.918 18.281 ;
 END
 END vccdgt_1p0.gds1022
 PIN vccdgt_1p0.gds1023
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.074 18.3635 6.114 18.5635 ;
 END
 END vccdgt_1p0.gds1023
 PIN vccdgt_1p0.gds1024
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.306 18.081 5.346 18.281 ;
 END
 END vccdgt_1p0.gds1024
 PIN vccdgt_1p0.gds1025
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.818 18.592 5.858 18.792 ;
 END
 END vccdgt_1p0.gds1025
 PIN vccdgt_1p0.gds1026
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.498 19.62 5.538 19.82 ;
 END
 END vccdgt_1p0.gds1026
 PIN vccdgt_1p0.gds1027
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.458 17.051 6.498 17.251 ;
 END
 END vccdgt_1p0.gds1027
 PIN vccdgt_1p0.gds1028
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.202 18.0345 6.242 18.2345 ;
 END
 END vccdgt_1p0.gds1028
 PIN vccdgt_1p0.gds1029
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.67 18.4455 6.71 18.6455 ;
 END
 END vccdgt_1p0.gds1029
 PIN vccdgt_1p0.gds1030
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 9.884 18.127 9.94 18.327 ;
 RECT 9.716 18.127 9.772 18.327 ;
 RECT 10.22 18.127 10.276 18.327 ;
 RECT 10.052 18.127 10.108 18.327 ;
 RECT 9.212 18.127 9.268 18.327 ;
 RECT 9.044 18.127 9.1 18.327 ;
 RECT 9.548 18.127 9.604 18.327 ;
 RECT 9.38 18.127 9.436 18.327 ;
 RECT 8.54 18.127 8.596 18.327 ;
 RECT 8.372 18.127 8.428 18.327 ;
 RECT 8.876 18.127 8.932 18.327 ;
 RECT 8.708 18.127 8.764 18.327 ;
 RECT 7.868 18.127 7.924 18.327 ;
 RECT 7.7 18.127 7.756 18.327 ;
 RECT 8.204 18.127 8.26 18.327 ;
 RECT 9.968 16.433 10.024 16.633 ;
 RECT 9.8 16.433 9.856 16.633 ;
 RECT 10.136 16.433 10.192 16.633 ;
 RECT 9.296 16.433 9.352 16.633 ;
 RECT 9.128 16.433 9.184 16.633 ;
 RECT 9.632 16.433 9.688 16.633 ;
 RECT 9.464 16.433 9.52 16.633 ;
 RECT 8.624 16.433 8.68 16.633 ;
 RECT 8.456 16.433 8.512 16.633 ;
 RECT 8.96 16.433 9.016 16.633 ;
 RECT 8.792 16.433 8.848 16.633 ;
 RECT 7.952 16.433 8.008 16.633 ;
 RECT 7.784 16.433 7.84 16.633 ;
 RECT 8.288 16.433 8.344 16.633 ;
 RECT 8.12 16.433 8.176 16.633 ;
 RECT 7.28 16.433 7.336 16.633 ;
 RECT 7.112 16.433 7.168 16.633 ;
 RECT 6.944 16.433 7 16.633 ;
 RECT 7.616 16.433 7.672 16.633 ;
 RECT 7.448 16.433 7.504 16.633 ;
 RECT 9.968 17.2925 10.024 17.4925 ;
 RECT 9.8 17.2915 9.856 17.4915 ;
 RECT 10.136 17.2925 10.192 17.4925 ;
 RECT 9.296 17.2925 9.352 17.4925 ;
 RECT 9.128 17.2915 9.184 17.4915 ;
 RECT 9.632 17.106 9.688 17.306 ;
 RECT 9.464 17.2925 9.52 17.4925 ;
 RECT 8.624 17.2925 8.68 17.4925 ;
 RECT 8.456 17.2915 8.512 17.4915 ;
 RECT 8.96 17.106 9.016 17.306 ;
 RECT 8.792 17.2925 8.848 17.4925 ;
 RECT 7.952 17.2925 8.008 17.4925 ;
 RECT 7.784 17.2915 7.84 17.4915 ;
 RECT 8.288 17.106 8.344 17.306 ;
 RECT 8.12 17.2925 8.176 17.4925 ;
 RECT 7.28 17.2925 7.336 17.4925 ;
 RECT 6.944 17.106 7 17.306 ;
 RECT 7.616 17.106 7.672 17.306 ;
 RECT 7.112 17.2915 7.168 17.4915 ;
 RECT 7.448 17.2925 7.504 17.4925 ;
 RECT 6.02 19.1975 6.076 19.3975 ;
 RECT 5.348 19.2485 5.404 19.4485 ;
 RECT 5.684 19.2765 5.74 19.4765 ;
 RECT 6.356 19.2765 6.412 19.4765 ;
 RECT 5.936 16.574 5.992 16.774 ;
 RECT 5.768 16.574 5.824 16.774 ;
 RECT 5.6 16.574 5.656 16.774 ;
 RECT 5.432 16.574 5.488 16.774 ;
 RECT 6.272 16.574 6.328 16.774 ;
 RECT 6.104 16.574 6.16 16.774 ;
 RECT 6.44 16.574 6.496 16.774 ;
 RECT 5.936 17.918 5.992 18.118 ;
 RECT 5.768 17.918 5.824 18.118 ;
 RECT 5.6 17.918 5.656 18.118 ;
 RECT 5.432 17.918 5.488 18.118 ;
 RECT 6.272 17.918 6.328 18.118 ;
 RECT 6.104 17.918 6.16 18.118 ;
 RECT 6.44 18.058 6.496 18.258 ;
 RECT 8.036 18.127 8.092 18.327 ;
 RECT 7.196 18.127 7.252 18.327 ;
 RECT 7.028 18.127 7.084 18.327 ;
 RECT 7.364 18.127 7.42 18.327 ;
 RECT 7.532 18.127 7.588 18.327 ;
 END
 END vccdgt_1p0.gds1030
 PIN vccdgt_1p0.gds1031
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.762 15.447 13.818 15.647 ;
 END
 END vccdgt_1p0.gds1031
 PIN vccdgt_1p0.gds1032
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.522 17.2285 14.578 17.4285 ;
 END
 END vccdgt_1p0.gds1032
 PIN vccdgt_1p0.gds1033
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.73 15.679 11.77 15.879 ;
 END
 END vccdgt_1p0.gds1033
 PIN vccdgt_1p0.gds1034
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.058 15.679 11.098 15.879 ;
 END
 END vccdgt_1p0.gds1034
 PIN vccdgt_1p0.gds1035
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.386 15.679 10.426 15.879 ;
 END
 END vccdgt_1p0.gds1035
 PIN vccdgt_1p0.gds1036
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.342 18.348 13.398 18.548 ;
 END
 END vccdgt_1p0.gds1036
 PIN vccdgt_1p0.gds1037
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.186 18.7195 15.226 18.9195 ;
 END
 END vccdgt_1p0.gds1037
 PIN vccdgt_1p0.gds1038
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.182 18.2595 14.238 18.4595 ;
 END
 END vccdgt_1p0.gds1038
 PIN vccdgt_1p0.gds1039
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.502 18.5525 13.558 18.7525 ;
 END
 END vccdgt_1p0.gds1039
 PIN vccdgt_1p0.gds1040
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.162 18.266 13.238 18.466 ;
 END
 END vccdgt_1p0.gds1040
 PIN vccdgt_1p0.gds1041
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.766 17.3945 14.806 17.5945 ;
 END
 END vccdgt_1p0.gds1041
 PIN vccdgt_1p0.gds1042
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.002 18.154 14.078 18.354 ;
 END
 END vccdgt_1p0.gds1042
 PIN vccdgt_1p0.gds1043
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.958 18.084 14.998 18.284 ;
 END
 END vccdgt_1p0.gds1043
 PIN vccdgt_1p0.gds1044
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.982 17.5555 12.042 17.7555 ;
 END
 END vccdgt_1p0.gds1044
 PIN vccdgt_1p0.gds1045
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.31 17.5555 11.37 17.7555 ;
 END
 END vccdgt_1p0.gds1045
 PIN vccdgt_1p0.gds1046
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.638 17.5555 10.698 17.7555 ;
 END
 END vccdgt_1p0.gds1046
 PIN vccdgt_1p0.gds1047
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.678 18.3175 12.718 18.5175 ;
 END
 END vccdgt_1p0.gds1047
 PIN vccdgt_1p0.gds1048
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.402 18.4715 12.462 18.6715 ;
 END
 END vccdgt_1p0.gds1048
 PIN vccdgt_1p0.gds1049
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 11.9 18.127 11.956 18.327 ;
 RECT 11.732 18.127 11.788 18.327 ;
 RECT 12.236 18.127 12.292 18.327 ;
 RECT 12.068 18.127 12.124 18.327 ;
 RECT 11.228 18.127 11.284 18.327 ;
 RECT 11.06 18.127 11.116 18.327 ;
 RECT 11.564 18.127 11.62 18.327 ;
 RECT 11.396 18.127 11.452 18.327 ;
 RECT 10.556 18.127 10.612 18.327 ;
 RECT 10.388 18.127 10.444 18.327 ;
 RECT 10.892 18.127 10.948 18.327 ;
 RECT 10.724 18.127 10.78 18.327 ;
 RECT 13.664 16.434 13.72 16.634 ;
 RECT 12.824 16.434 12.88 16.634 ;
 RECT 13.496 16.434 13.552 16.634 ;
 RECT 13.16 16.434 13.216 16.634 ;
 RECT 12.992 16.434 13.048 16.634 ;
 RECT 14.168 16.434 14.224 16.634 ;
 RECT 14 16.434 14.056 16.634 ;
 RECT 15.176 16.434 15.232 16.634 ;
 RECT 15.008 16.434 15.064 16.634 ;
 RECT 14.84 16.434 14.896 16.634 ;
 RECT 14.672 16.431 14.728 16.631 ;
 RECT 14.504 16.434 14.56 16.634 ;
 RECT 11.984 16.433 12.04 16.633 ;
 RECT 11.816 16.433 11.872 16.633 ;
 RECT 12.32 16.433 12.376 16.633 ;
 RECT 12.152 16.433 12.208 16.633 ;
 RECT 11.312 16.433 11.368 16.633 ;
 RECT 11.144 16.433 11.2 16.633 ;
 RECT 11.648 16.433 11.704 16.633 ;
 RECT 11.48 16.433 11.536 16.633 ;
 RECT 10.64 16.433 10.696 16.633 ;
 RECT 10.472 16.433 10.528 16.633 ;
 RECT 10.976 16.433 11.032 16.633 ;
 RECT 10.808 16.433 10.864 16.633 ;
 RECT 10.304 16.433 10.36 16.633 ;
 RECT 13.664 17.63 13.72 17.83 ;
 RECT 12.824 17.63 12.88 17.83 ;
 RECT 14.336 17.742 14.392 17.942 ;
 RECT 14.672 17.6715 14.728 17.8715 ;
 RECT 12.488 17.3055 12.544 17.5055 ;
 RECT 12.656 17.533 12.712 17.733 ;
 RECT 14 19.04 14.056 19.24 ;
 RECT 14.756 20.417 14.812 20.617 ;
 RECT 14.924 19.984 14.98 20.184 ;
 RECT 14 20.3 14.056 20.5 ;
 RECT 14.588 20.417 14.644 20.617 ;
 RECT 14.42 20.404 14.476 20.604 ;
 RECT 14.756 19.157 14.812 19.357 ;
 RECT 14.924 18.724 14.98 18.924 ;
 RECT 14.588 19.157 14.644 19.357 ;
 RECT 14.42 19.144 14.476 19.344 ;
 RECT 12.404 16.183 12.46 16.383 ;
 RECT 13.328 16.63 13.384 16.83 ;
 RECT 14.168 17.6435 14.224 17.8435 ;
 RECT 14 17.5755 14.056 17.7755 ;
 RECT 13.832 17.472 13.888 17.672 ;
 RECT 14.84 17.533 14.896 17.733 ;
 RECT 14.504 17.5895 14.56 17.7895 ;
 RECT 15.008 17.533 15.064 17.733 ;
 RECT 15.176 17.5895 15.232 17.7895 ;
 RECT 11.984 17.2925 12.04 17.4925 ;
 RECT 11.816 17.2915 11.872 17.4915 ;
 RECT 12.32 17.106 12.376 17.306 ;
 RECT 12.152 17.2925 12.208 17.4925 ;
 RECT 11.312 17.2925 11.368 17.4925 ;
 RECT 11.144 17.2915 11.2 17.4915 ;
 RECT 11.648 17.106 11.704 17.306 ;
 RECT 11.48 17.2925 11.536 17.4925 ;
 RECT 10.64 17.2925 10.696 17.4925 ;
 RECT 10.472 17.2915 10.528 17.4915 ;
 RECT 10.976 17.106 11.032 17.306 ;
 RECT 10.808 17.2925 10.864 17.4925 ;
 RECT 10.304 17.106 10.36 17.306 ;
 END
 END vccdgt_1p0.gds1049
 PIN vccdgt_1p0.gds1050
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.626 15.679 19.666 15.879 ;
 END
 END vccdgt_1p0.gds1050
 PIN vccdgt_1p0.gds1051
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 19.666 16.57 19.866 ;
 END
 END vccdgt_1p0.gds1051
 PIN vccdgt_1p0.gds1052
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.866 18.185 15.926 18.385 ;
 END
 END vccdgt_1p0.gds1052
 PIN vccdgt_1p0.gds1053
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.954 15.679 18.994 15.879 ;
 END
 END vccdgt_1p0.gds1053
 PIN vccdgt_1p0.gds1054
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.282 15.679 18.322 15.879 ;
 END
 END vccdgt_1p0.gds1054
 PIN vccdgt_1p0.gds1055
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.838 19.5775 16.894 19.7775 ;
 END
 END vccdgt_1p0.gds1055
 PIN vccdgt_1p0.gds1056
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.674 18.911 16.734 19.111 ;
 END
 END vccdgt_1p0.gds1056
 PIN vccdgt_1p0.gds1057
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.018 19.3865 17.074 19.5865 ;
 END
 END vccdgt_1p0.gds1057
 PIN vccdgt_1p0.gds1058
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.878 17.5555 19.938 17.7555 ;
 END
 END vccdgt_1p0.gds1058
 PIN vccdgt_1p0.gds1059
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 17.697 16.57 17.897 ;
 END
 END vccdgt_1p0.gds1059
 PIN vccdgt_1p0.gds1060
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.03 17.965 16.076 18.165 ;
 END
 END vccdgt_1p0.gds1060
 PIN vccdgt_1p0.gds1061
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.314 17.6915 15.354 17.8915 ;
 END
 END vccdgt_1p0.gds1061
 PIN vccdgt_1p0.gds1062
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.338 18.1605 17.414 18.3605 ;
 END
 END vccdgt_1p0.gds1062
 PIN vccdgt_1p0.gds1063
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.114 18.2535 18.174 18.4535 ;
 END
 END vccdgt_1p0.gds1063
 PIN vccdgt_1p0.gds1064
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.858 19.4835 17.898 19.6835 ;
 END
 END vccdgt_1p0.gds1064
 PIN vccdgt_1p0.gds1065
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.522 17.757 15.582 17.957 ;
 END
 END vccdgt_1p0.gds1065
 PIN vccdgt_1p0.gds1066
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.598 17.845 17.654 18.045 ;
 END
 END vccdgt_1p0.gds1066
 PIN vccdgt_1p0.gds1067
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.178 17.8845 17.234 18.0845 ;
 END
 END vccdgt_1p0.gds1067
 PIN vccdgt_1p0.gds1068
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.206 17.5555 19.266 17.7555 ;
 END
 END vccdgt_1p0.gds1068
 PIN vccdgt_1p0.gds1069
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.534 17.5555 18.594 17.7555 ;
 END
 END vccdgt_1p0.gds1069
 PIN vccdgt_1p0.gds1070
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 19.796 18.127 19.852 18.327 ;
 RECT 19.628 18.127 19.684 18.327 ;
 RECT 19.964 18.127 20.02 18.327 ;
 RECT 20.132 18.127 20.188 18.327 ;
 RECT 19.124 18.127 19.18 18.327 ;
 RECT 18.956 18.127 19.012 18.327 ;
 RECT 19.292 18.127 19.348 18.327 ;
 RECT 19.46 18.127 19.516 18.327 ;
 RECT 18.452 18.127 18.508 18.327 ;
 RECT 18.284 18.127 18.34 18.327 ;
 RECT 18.788 18.127 18.844 18.327 ;
 RECT 18.62 18.127 18.676 18.327 ;
 RECT 19.88 16.433 19.936 16.633 ;
 RECT 19.712 16.433 19.768 16.633 ;
 RECT 20.216 16.433 20.272 16.633 ;
 RECT 20.048 16.433 20.104 16.633 ;
 RECT 16.1 16.434 16.156 16.634 ;
 RECT 15.764 16.434 15.82 16.634 ;
 RECT 15.596 16.434 15.652 16.634 ;
 RECT 15.428 16.434 15.484 16.634 ;
 RECT 16.772 16.434 16.828 16.634 ;
 RECT 16.604 16.434 16.66 16.634 ;
 RECT 16.436 16.434 16.492 16.634 ;
 RECT 16.268 16.434 16.324 16.634 ;
 RECT 17.276 16.471 17.332 16.653 ;
 RECT 17.024 16.471 17.08 16.653 ;
 RECT 17.612 16.435 17.668 16.635 ;
 RECT 19.208 16.433 19.264 16.633 ;
 RECT 19.04 16.433 19.096 16.633 ;
 RECT 19.544 16.433 19.6 16.633 ;
 RECT 19.376 16.433 19.432 16.633 ;
 RECT 18.536 16.433 18.592 16.633 ;
 RECT 18.368 16.433 18.424 16.633 ;
 RECT 18.2 16.433 18.256 16.633 ;
 RECT 18.872 16.433 18.928 16.633 ;
 RECT 18.704 16.433 18.76 16.633 ;
 RECT 18.032 17.783 18.088 17.983 ;
 RECT 19.88 17.2925 19.936 17.4925 ;
 RECT 19.712 17.2915 19.768 17.4915 ;
 RECT 20.216 17.106 20.272 17.306 ;
 RECT 20.048 17.2925 20.104 17.4925 ;
 RECT 15.68 17.6715 15.736 17.8715 ;
 RECT 15.344 17.601 15.4 17.801 ;
 RECT 17.36 17.5645 17.416 17.7645 ;
 RECT 17.528 17.5645 17.584 17.7645 ;
 RECT 16.1 19.157 16.156 19.357 ;
 RECT 15.764 20.06 15.82 20.26 ;
 RECT 18.116 15.621 18.172 15.821 ;
 RECT 15.512 20.312 15.568 20.512 ;
 RECT 15.26 20.399 15.316 20.599 ;
 RECT 16.1 20.417 16.156 20.617 ;
 RECT 15.932 19.22 15.988 19.42 ;
 RECT 15.764 18.8 15.82 19 ;
 RECT 15.512 19.052 15.568 19.252 ;
 RECT 15.26 19.139 15.316 19.339 ;
 RECT 16.856 17.533 16.912 17.733 ;
 RECT 15.512 17.5895 15.568 17.7895 ;
 RECT 16.016 17.533 16.072 17.733 ;
 RECT 15.848 17.533 15.904 17.733 ;
 RECT 16.688 17.533 16.744 17.733 ;
 RECT 16.52 17.533 16.576 17.733 ;
 RECT 16.352 17.533 16.408 17.733 ;
 RECT 16.184 17.533 16.24 17.733 ;
 RECT 17.696 17.4855 17.752 17.6855 ;
 RECT 17.192 17.4855 17.248 17.6855 ;
 RECT 17.864 17.4855 17.92 17.6855 ;
 RECT 19.208 17.2925 19.264 17.4925 ;
 RECT 19.04 17.2915 19.096 17.4915 ;
 RECT 19.544 17.106 19.6 17.306 ;
 RECT 19.376 17.2925 19.432 17.4925 ;
 RECT 18.536 17.2925 18.592 17.4925 ;
 RECT 18.368 17.2915 18.424 17.4915 ;
 RECT 18.2 17.106 18.256 17.306 ;
 RECT 18.872 17.106 18.928 17.306 ;
 RECT 18.704 17.2925 18.76 17.4925 ;
 RECT 17.024 17.498 17.08 17.698 ;
 END
 END vccdgt_1p0.gds1070
 PIN vccdgt_1p0.gds1071
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.078 15.679 24.118 15.879 ;
 END
 END vccdgt_1p0.gds1071
 PIN vccdgt_1p0.gds1072
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.986 15.679 23.026 15.879 ;
 END
 END vccdgt_1p0.gds1072
 PIN vccdgt_1p0.gds1073
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.75 15.679 24.79 15.879 ;
 END
 END vccdgt_1p0.gds1073
 PIN vccdgt_1p0.gds1074
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.314 15.679 22.354 15.879 ;
 END
 END vccdgt_1p0.gds1074
 PIN vccdgt_1p0.gds1075
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.642 15.679 21.682 15.879 ;
 END
 END vccdgt_1p0.gds1075
 PIN vccdgt_1p0.gds1076
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.97 15.679 21.01 15.879 ;
 END
 END vccdgt_1p0.gds1076
 PIN vccdgt_1p0.gds1077
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.298 15.679 20.338 15.879 ;
 END
 END vccdgt_1p0.gds1077
 PIN vccdgt_1p0.gds1078
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.002 17.5555 25.062 17.7555 ;
 END
 END vccdgt_1p0.gds1078
 PIN vccdgt_1p0.gds1079
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.33 17.5555 24.39 17.7555 ;
 END
 END vccdgt_1p0.gds1079
 PIN vccdgt_1p0.gds1080
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.238 17.5555 23.298 17.7555 ;
 END
 END vccdgt_1p0.gds1080
 PIN vccdgt_1p0.gds1081
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.566 17.5555 22.626 17.7555 ;
 END
 END vccdgt_1p0.gds1081
 PIN vccdgt_1p0.gds1082
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.894 17.5555 21.954 17.7555 ;
 END
 END vccdgt_1p0.gds1082
 PIN vccdgt_1p0.gds1083
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.222 17.5555 21.282 17.7555 ;
 END
 END vccdgt_1p0.gds1083
 PIN vccdgt_1p0.gds1084
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.55 17.5555 20.61 17.7555 ;
 END
 END vccdgt_1p0.gds1084
 PIN vccdgt_1p0.gds1085
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.93 18.16 23.97 18.36 ;
 END
 END vccdgt_1p0.gds1085
 PIN vccdgt_1p0.gds1086
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.658 17.915 23.698 18.115 ;
 END
 END vccdgt_1p0.gds1086
 PIN vccdgt_1p0.gds1087
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 24.92 18.127 24.976 18.327 ;
 RECT 24.752 18.127 24.808 18.327 ;
 RECT 25.088 18.127 25.144 18.327 ;
 RECT 24.248 18.127 24.304 18.327 ;
 RECT 24.08 18.127 24.136 18.327 ;
 RECT 24.416 18.127 24.472 18.327 ;
 RECT 24.584 18.127 24.64 18.327 ;
 RECT 23.156 18.127 23.212 18.327 ;
 RECT 22.988 18.127 23.044 18.327 ;
 RECT 23.324 18.127 23.38 18.327 ;
 RECT 23.492 18.127 23.548 18.327 ;
 RECT 22.484 18.127 22.54 18.327 ;
 RECT 22.316 18.127 22.372 18.327 ;
 RECT 22.652 18.127 22.708 18.327 ;
 RECT 22.82 18.127 22.876 18.327 ;
 RECT 21.812 18.127 21.868 18.327 ;
 RECT 21.644 18.127 21.7 18.327 ;
 RECT 21.98 18.127 22.036 18.327 ;
 RECT 22.148 18.127 22.204 18.327 ;
 RECT 21.14 18.127 21.196 18.327 ;
 RECT 20.972 18.127 21.028 18.327 ;
 RECT 21.308 18.127 21.364 18.327 ;
 RECT 21.476 18.127 21.532 18.327 ;
 RECT 20.468 18.127 20.524 18.327 ;
 RECT 20.636 18.127 20.692 18.327 ;
 RECT 20.804 18.127 20.86 18.327 ;
 RECT 20.3 18.127 20.356 18.327 ;
 RECT 25.004 16.433 25.06 16.633 ;
 RECT 24.836 16.433 24.892 16.633 ;
 RECT 25.172 16.433 25.228 16.633 ;
 RECT 24.332 16.433 24.388 16.633 ;
 RECT 24.164 16.433 24.22 16.633 ;
 RECT 23.996 16.433 24.052 16.633 ;
 RECT 24.668 16.433 24.724 16.633 ;
 RECT 24.5 16.433 24.556 16.633 ;
 RECT 23.24 16.433 23.296 16.633 ;
 RECT 23.072 16.433 23.128 16.633 ;
 RECT 23.576 16.433 23.632 16.633 ;
 RECT 23.408 16.433 23.464 16.633 ;
 RECT 22.568 16.433 22.624 16.633 ;
 RECT 22.4 16.433 22.456 16.633 ;
 RECT 22.904 16.433 22.96 16.633 ;
 RECT 22.736 16.433 22.792 16.633 ;
 RECT 21.896 16.433 21.952 16.633 ;
 RECT 21.728 16.433 21.784 16.633 ;
 RECT 22.232 16.433 22.288 16.633 ;
 RECT 22.064 16.433 22.12 16.633 ;
 RECT 21.224 16.433 21.28 16.633 ;
 RECT 21.056 16.433 21.112 16.633 ;
 RECT 21.56 16.433 21.616 16.633 ;
 RECT 21.392 16.433 21.448 16.633 ;
 RECT 20.552 16.433 20.608 16.633 ;
 RECT 20.888 16.433 20.944 16.633 ;
 RECT 20.72 16.433 20.776 16.633 ;
 RECT 20.384 16.433 20.44 16.633 ;
 RECT 25.004 17.2925 25.06 17.4925 ;
 RECT 24.836 17.2915 24.892 17.4915 ;
 RECT 25.172 17.2925 25.228 17.4925 ;
 RECT 24.332 17.2925 24.388 17.4925 ;
 RECT 24.164 17.2915 24.22 17.4915 ;
 RECT 23.996 17.106 24.052 17.306 ;
 RECT 24.668 17.106 24.724 17.306 ;
 RECT 24.5 17.2925 24.556 17.4925 ;
 RECT 23.24 17.2925 23.296 17.4925 ;
 RECT 23.072 17.2915 23.128 17.4915 ;
 RECT 23.576 17.106 23.632 17.306 ;
 RECT 23.408 17.2925 23.464 17.4925 ;
 RECT 22.568 17.2925 22.624 17.4925 ;
 RECT 22.4 17.2915 22.456 17.4915 ;
 RECT 22.904 17.106 22.96 17.306 ;
 RECT 22.736 17.2925 22.792 17.4925 ;
 RECT 21.896 17.2925 21.952 17.4925 ;
 RECT 21.728 17.2915 21.784 17.4915 ;
 RECT 22.232 17.106 22.288 17.306 ;
 RECT 22.064 17.2925 22.12 17.4925 ;
 RECT 21.224 17.2925 21.28 17.4925 ;
 RECT 21.056 17.2915 21.112 17.4915 ;
 RECT 21.56 17.106 21.616 17.306 ;
 RECT 21.392 17.2925 21.448 17.4925 ;
 RECT 20.552 17.2925 20.608 17.4925 ;
 RECT 20.888 17.106 20.944 17.306 ;
 RECT 20.72 17.2925 20.776 17.4925 ;
 RECT 20.384 17.2915 20.44 17.4915 ;
 RECT 23.828 16.434 23.884 16.634 ;
 RECT 23.912 17.2105 23.968 17.4105 ;
 RECT 23.66 17.3245 23.716 17.5245 ;
 END
 END vccdgt_1p0.gds1087
 PIN vccdgt_1p0.gds1088
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.782 15.679 28.822 15.879 ;
 END
 END vccdgt_1p0.gds1088
 PIN vccdgt_1p0.gds1089
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.11 15.679 28.15 15.879 ;
 END
 END vccdgt_1p0.gds1089
 PIN vccdgt_1p0.gds1090
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.438 15.679 27.478 15.879 ;
 END
 END vccdgt_1p0.gds1090
 PIN vccdgt_1p0.gds1091
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.766 15.679 26.806 15.879 ;
 END
 END vccdgt_1p0.gds1091
 PIN vccdgt_1p0.gds1092
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.094 15.679 26.134 15.879 ;
 END
 END vccdgt_1p0.gds1092
 PIN vccdgt_1p0.gds1093
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.422 15.679 25.462 15.879 ;
 END
 END vccdgt_1p0.gds1093
 PIN vccdgt_1p0.gds1094
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.034 17.5555 29.094 17.7555 ;
 END
 END vccdgt_1p0.gds1094
 PIN vccdgt_1p0.gds1095
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.362 17.5555 28.422 17.7555 ;
 END
 END vccdgt_1p0.gds1095
 PIN vccdgt_1p0.gds1096
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.69 17.5555 27.75 17.7555 ;
 END
 END vccdgt_1p0.gds1096
 PIN vccdgt_1p0.gds1097
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.018 17.5555 27.078 17.7555 ;
 END
 END vccdgt_1p0.gds1097
 PIN vccdgt_1p0.gds1098
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.346 17.5555 26.406 17.7555 ;
 END
 END vccdgt_1p0.gds1098
 PIN vccdgt_1p0.gds1099
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.674 17.5555 25.734 17.7555 ;
 END
 END vccdgt_1p0.gds1099
 PIN vccdgt_1p0.gds1100
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.214 18.266 30.29 18.466 ;
 END
 END vccdgt_1p0.gds1100
 PIN vccdgt_1p0.gds1101
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.73 18.3175 29.77 18.5175 ;
 END
 END vccdgt_1p0.gds1101
 PIN vccdgt_1p0.gds1102
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.454 18.4715 29.514 18.6715 ;
 END
 END vccdgt_1p0.gds1102
 PIN vccdgt_1p0.gds1103
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 28.952 18.127 29.008 18.327 ;
 RECT 28.784 18.127 28.84 18.327 ;
 RECT 29.12 18.127 29.176 18.327 ;
 RECT 29.288 18.127 29.344 18.327 ;
 RECT 28.28 18.127 28.336 18.327 ;
 RECT 28.112 18.127 28.168 18.327 ;
 RECT 28.448 18.127 28.504 18.327 ;
 RECT 28.616 18.127 28.672 18.327 ;
 RECT 27.608 18.127 27.664 18.327 ;
 RECT 27.44 18.127 27.496 18.327 ;
 RECT 27.776 18.127 27.832 18.327 ;
 RECT 27.944 18.127 28 18.327 ;
 RECT 26.936 18.127 26.992 18.327 ;
 RECT 26.768 18.127 26.824 18.327 ;
 RECT 27.104 18.127 27.16 18.327 ;
 RECT 27.272 18.127 27.328 18.327 ;
 RECT 26.264 18.127 26.32 18.327 ;
 RECT 26.096 18.127 26.152 18.327 ;
 RECT 26.432 18.127 26.488 18.327 ;
 RECT 26.6 18.127 26.656 18.327 ;
 RECT 25.592 18.127 25.648 18.327 ;
 RECT 25.424 18.127 25.48 18.327 ;
 RECT 25.76 18.127 25.816 18.327 ;
 RECT 25.928 18.127 25.984 18.327 ;
 RECT 25.256 18.127 25.312 18.327 ;
 RECT 29.876 16.434 29.932 16.634 ;
 RECT 30.212 16.434 30.268 16.634 ;
 RECT 30.044 16.434 30.1 16.634 ;
 RECT 29.036 16.433 29.092 16.633 ;
 RECT 28.868 16.433 28.924 16.633 ;
 RECT 29.372 16.433 29.428 16.633 ;
 RECT 29.204 16.433 29.26 16.633 ;
 RECT 28.364 16.433 28.42 16.633 ;
 RECT 28.196 16.433 28.252 16.633 ;
 RECT 28.7 16.433 28.756 16.633 ;
 RECT 28.532 16.433 28.588 16.633 ;
 RECT 27.692 16.433 27.748 16.633 ;
 RECT 27.524 16.433 27.58 16.633 ;
 RECT 28.028 16.433 28.084 16.633 ;
 RECT 27.86 16.433 27.916 16.633 ;
 RECT 27.02 16.433 27.076 16.633 ;
 RECT 26.852 16.433 26.908 16.633 ;
 RECT 27.356 16.433 27.412 16.633 ;
 RECT 27.188 16.433 27.244 16.633 ;
 RECT 26.348 16.433 26.404 16.633 ;
 RECT 26.18 16.433 26.236 16.633 ;
 RECT 26.684 16.433 26.74 16.633 ;
 RECT 26.516 16.433 26.572 16.633 ;
 RECT 25.676 16.433 25.732 16.633 ;
 RECT 25.508 16.433 25.564 16.633 ;
 RECT 26.012 16.433 26.068 16.633 ;
 RECT 25.844 16.433 25.9 16.633 ;
 RECT 25.34 16.433 25.396 16.633 ;
 RECT 29.876 17.63 29.932 17.83 ;
 RECT 29.036 17.2925 29.092 17.4925 ;
 RECT 28.868 17.2915 28.924 17.4915 ;
 RECT 29.372 17.106 29.428 17.306 ;
 RECT 29.204 17.2925 29.26 17.4925 ;
 RECT 28.364 17.2925 28.42 17.4925 ;
 RECT 28.196 17.2915 28.252 17.4915 ;
 RECT 28.7 17.106 28.756 17.306 ;
 RECT 28.532 17.2925 28.588 17.4925 ;
 RECT 27.692 17.2925 27.748 17.4925 ;
 RECT 27.524 17.2915 27.58 17.4915 ;
 RECT 28.028 17.106 28.084 17.306 ;
 RECT 27.86 17.2925 27.916 17.4925 ;
 RECT 27.02 17.2925 27.076 17.4925 ;
 RECT 26.852 17.2915 26.908 17.4915 ;
 RECT 27.356 17.106 27.412 17.306 ;
 RECT 27.188 17.2925 27.244 17.4925 ;
 RECT 26.348 17.2925 26.404 17.4925 ;
 RECT 26.18 17.2915 26.236 17.4915 ;
 RECT 26.684 17.106 26.74 17.306 ;
 RECT 26.516 17.2925 26.572 17.4925 ;
 RECT 25.676 17.2925 25.732 17.4925 ;
 RECT 25.508 17.2915 25.564 17.4915 ;
 RECT 26.012 17.106 26.068 17.306 ;
 RECT 25.844 17.2925 25.9 17.4925 ;
 RECT 25.34 17.106 25.396 17.306 ;
 RECT 29.54 17.3055 29.596 17.5055 ;
 RECT 29.708 17.533 29.764 17.733 ;
 RECT 29.456 16.183 29.512 16.383 ;
 END
 END vccdgt_1p0.gds1103
 PIN vccdgt_1p0.gds1104
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.814 15.447 30.87 15.647 ;
 END
 END vccdgt_1p0.gds1104
 PIN vccdgt_1p0.gds1105
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 19.666 33.622 19.866 ;
 END
 END vccdgt_1p0.gds1105
 PIN vccdgt_1p0.gds1106
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.574 17.2285 31.63 17.4285 ;
 END
 END vccdgt_1p0.gds1106
 PIN vccdgt_1p0.gds1107
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.918 18.185 32.978 18.385 ;
 END
 END vccdgt_1p0.gds1107
 PIN vccdgt_1p0.gds1108
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.238 18.664 32.278 18.864 ;
 END
 END vccdgt_1p0.gds1108
 PIN vccdgt_1p0.gds1109
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.394 18.348 30.45 18.548 ;
 END
 END vccdgt_1p0.gds1109
 PIN vccdgt_1p0.gds1110
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.89 19.5775 33.946 19.7775 ;
 END
 END vccdgt_1p0.gds1110
 PIN vccdgt_1p0.gds1111
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.726 18.911 33.786 19.111 ;
 END
 END vccdgt_1p0.gds1111
 PIN vccdgt_1p0.gds1112
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.07 19.3865 34.126 19.5865 ;
 END
 END vccdgt_1p0.gds1112
 PIN vccdgt_1p0.gds1113
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 17.697 33.622 17.897 ;
 END
 END vccdgt_1p0.gds1113
 PIN vccdgt_1p0.gds1114
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.39 18.1605 34.466 18.3605 ;
 END
 END vccdgt_1p0.gds1114
 PIN vccdgt_1p0.gds1115
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.082 17.965 33.128 18.165 ;
 END
 END vccdgt_1p0.gds1115
 PIN vccdgt_1p0.gds1116
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.366 18.5935 32.406 18.7935 ;
 END
 END vccdgt_1p0.gds1116
 PIN vccdgt_1p0.gds1117
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.554 18.5525 30.61 18.7525 ;
 END
 END vccdgt_1p0.gds1117
 PIN vccdgt_1p0.gds1118
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.818 17.3945 31.858 17.5945 ;
 END
 END vccdgt_1p0.gds1118
 PIN vccdgt_1p0.gds1119
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.234 18.2595 31.29 18.4595 ;
 END
 END vccdgt_1p0.gds1119
 PIN vccdgt_1p0.gds1120
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.91 19.4835 34.95 19.6835 ;
 END
 END vccdgt_1p0.gds1120
 PIN vccdgt_1p0.gds1121
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.574 17.757 32.634 17.957 ;
 END
 END vccdgt_1p0.gds1121
 PIN vccdgt_1p0.gds1122
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.65 17.845 34.706 18.045 ;
 END
 END vccdgt_1p0.gds1122
 PIN vccdgt_1p0.gds1123
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.01 18.084 32.05 18.284 ;
 END
 END vccdgt_1p0.gds1123
 PIN vccdgt_1p0.gds1124
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.166 18.2535 35.226 18.4535 ;
 END
 END vccdgt_1p0.gds1124
 PIN vccdgt_1p0.gds1125
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.054 18.154 31.13 18.354 ;
 END
 END vccdgt_1p0.gds1125
 PIN vccdgt_1p0.gds1126
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.23 17.8845 34.286 18.0845 ;
 END
 END vccdgt_1p0.gds1126
 PIN vccdgt_1p0.gds1127
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 30.716 16.434 30.772 16.634 ;
 RECT 30.548 16.434 30.604 16.634 ;
 RECT 31.22 16.434 31.276 16.634 ;
 RECT 31.052 16.434 31.108 16.634 ;
 RECT 32.228 16.434 32.284 16.634 ;
 RECT 32.06 16.434 32.116 16.634 ;
 RECT 31.892 16.434 31.948 16.634 ;
 RECT 31.724 16.431 31.78 16.631 ;
 RECT 31.556 16.434 31.612 16.634 ;
 RECT 33.152 16.434 33.208 16.634 ;
 RECT 32.816 16.434 32.872 16.634 ;
 RECT 32.648 16.434 32.704 16.634 ;
 RECT 32.48 16.434 32.536 16.634 ;
 RECT 33.824 16.434 33.88 16.634 ;
 RECT 33.656 16.434 33.712 16.634 ;
 RECT 33.488 16.434 33.544 16.634 ;
 RECT 33.32 16.434 33.376 16.634 ;
 RECT 34.328 16.471 34.384 16.653 ;
 RECT 34.076 16.471 34.132 16.653 ;
 RECT 34.664 16.435 34.72 16.635 ;
 RECT 30.716 17.63 30.772 17.83 ;
 RECT 31.388 17.742 31.444 17.942 ;
 RECT 35.084 17.783 35.14 17.983 ;
 RECT 31.22 17.6435 31.276 17.8435 ;
 RECT 31.052 17.5755 31.108 17.7755 ;
 RECT 30.884 17.472 30.94 17.672 ;
 RECT 33.152 19.157 33.208 19.357 ;
 RECT 31.052 19.04 31.108 19.24 ;
 RECT 31.976 19.984 32.032 20.184 ;
 RECT 32.816 20.06 32.872 20.26 ;
 RECT 31.052 20.3 31.108 20.5 ;
 RECT 31.808 20.417 31.864 20.617 ;
 RECT 33.152 20.417 33.208 20.617 ;
 RECT 31.64 20.417 31.696 20.617 ;
 RECT 31.472 20.404 31.528 20.604 ;
 RECT 32.564 20.312 32.62 20.512 ;
 RECT 32.312 20.399 32.368 20.599 ;
 RECT 31.808 19.157 31.864 19.357 ;
 RECT 32.984 19.22 33.04 19.42 ;
 RECT 31.976 18.724 32.032 18.924 ;
 RECT 32.816 18.8 32.872 19 ;
 RECT 32.564 19.052 32.62 19.252 ;
 RECT 32.312 19.139 32.368 19.339 ;
 RECT 31.64 19.157 31.696 19.357 ;
 RECT 31.472 19.144 31.528 19.344 ;
 RECT 35.168 15.621 35.224 15.821 ;
 RECT 31.892 17.533 31.948 17.733 ;
 RECT 31.556 17.5895 31.612 17.7895 ;
 RECT 31.724 17.6715 31.78 17.8715 ;
 RECT 32.06 17.533 32.116 17.733 ;
 RECT 32.228 17.5895 32.284 17.7895 ;
 RECT 33.908 17.533 33.964 17.733 ;
 RECT 32.732 17.6715 32.788 17.8715 ;
 RECT 32.396 17.601 32.452 17.801 ;
 RECT 32.564 17.5895 32.62 17.7895 ;
 RECT 33.068 17.533 33.124 17.733 ;
 RECT 32.9 17.533 32.956 17.733 ;
 RECT 33.74 17.533 33.796 17.733 ;
 RECT 33.572 17.533 33.628 17.733 ;
 RECT 33.404 17.533 33.46 17.733 ;
 RECT 33.236 17.533 33.292 17.733 ;
 RECT 34.748 17.4855 34.804 17.6855 ;
 RECT 34.412 17.5645 34.468 17.7645 ;
 RECT 34.076 17.498 34.132 17.698 ;
 RECT 34.58 17.5645 34.636 17.7645 ;
 RECT 34.244 17.4855 34.3 17.6855 ;
 RECT 34.916 17.4855 34.972 17.6855 ;
 RECT 30.38 16.63 30.436 16.83 ;
 END
 END vccdgt_1p0.gds1127
 PIN vccdgt_1p0.gds1128
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.366 15.679 39.406 15.879 ;
 END
 END vccdgt_1p0.gds1128
 PIN vccdgt_1p0.gds1129
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.694 15.679 38.734 15.879 ;
 END
 END vccdgt_1p0.gds1129
 PIN vccdgt_1p0.gds1130
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.022 15.679 38.062 15.879 ;
 END
 END vccdgt_1p0.gds1130
 PIN vccdgt_1p0.gds1131
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.35 15.679 37.39 15.879 ;
 END
 END vccdgt_1p0.gds1131
 PIN vccdgt_1p0.gds1132
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.678 15.679 36.718 15.879 ;
 END
 END vccdgt_1p0.gds1132
 PIN vccdgt_1p0.gds1133
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.006 15.679 36.046 15.879 ;
 END
 END vccdgt_1p0.gds1133
 PIN vccdgt_1p0.gds1134
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.038 15.679 40.078 15.879 ;
 END
 END vccdgt_1p0.gds1134
 PIN vccdgt_1p0.gds1135
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.334 15.679 35.374 15.879 ;
 END
 END vccdgt_1p0.gds1135
 PIN vccdgt_1p0.gds1136
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.618 17.5555 39.678 17.7555 ;
 END
 END vccdgt_1p0.gds1136
 PIN vccdgt_1p0.gds1137
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.946 17.5555 39.006 17.7555 ;
 END
 END vccdgt_1p0.gds1137
 PIN vccdgt_1p0.gds1138
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.274 17.5555 38.334 17.7555 ;
 END
 END vccdgt_1p0.gds1138
 PIN vccdgt_1p0.gds1139
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.602 17.5555 37.662 17.7555 ;
 END
 END vccdgt_1p0.gds1139
 PIN vccdgt_1p0.gds1140
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.93 17.5555 36.99 17.7555 ;
 END
 END vccdgt_1p0.gds1140
 PIN vccdgt_1p0.gds1141
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.258 17.5555 36.318 17.7555 ;
 END
 END vccdgt_1p0.gds1141
 PIN vccdgt_1p0.gds1142
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.586 17.5555 35.646 17.7555 ;
 END
 END vccdgt_1p0.gds1142
 PIN vccdgt_1p0.gds1143
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 40.208 18.127 40.264 18.327 ;
 RECT 40.04 18.127 40.096 18.327 ;
 RECT 39.536 18.127 39.592 18.327 ;
 RECT 39.368 18.127 39.424 18.327 ;
 RECT 39.704 18.127 39.76 18.327 ;
 RECT 39.872 18.127 39.928 18.327 ;
 RECT 38.864 18.127 38.92 18.327 ;
 RECT 38.696 18.127 38.752 18.327 ;
 RECT 39.032 18.127 39.088 18.327 ;
 RECT 39.2 18.127 39.256 18.327 ;
 RECT 38.192 18.127 38.248 18.327 ;
 RECT 38.024 18.127 38.08 18.327 ;
 RECT 38.36 18.127 38.416 18.327 ;
 RECT 38.528 18.127 38.584 18.327 ;
 RECT 37.52 18.127 37.576 18.327 ;
 RECT 37.352 18.127 37.408 18.327 ;
 RECT 37.688 18.127 37.744 18.327 ;
 RECT 37.856 18.127 37.912 18.327 ;
 RECT 36.848 18.127 36.904 18.327 ;
 RECT 36.68 18.127 36.736 18.327 ;
 RECT 37.016 18.127 37.072 18.327 ;
 RECT 37.184 18.127 37.24 18.327 ;
 RECT 36.176 18.127 36.232 18.327 ;
 RECT 36.008 18.127 36.064 18.327 ;
 RECT 36.344 18.127 36.4 18.327 ;
 RECT 36.512 18.127 36.568 18.327 ;
 RECT 35.504 18.127 35.56 18.327 ;
 RECT 35.336 18.127 35.392 18.327 ;
 RECT 35.84 18.127 35.896 18.327 ;
 RECT 35.672 18.127 35.728 18.327 ;
 RECT 40.124 16.433 40.18 16.633 ;
 RECT 39.62 16.433 39.676 16.633 ;
 RECT 39.452 16.433 39.508 16.633 ;
 RECT 39.956 16.433 40.012 16.633 ;
 RECT 39.788 16.433 39.844 16.633 ;
 RECT 38.948 16.433 39.004 16.633 ;
 RECT 38.78 16.433 38.836 16.633 ;
 RECT 39.284 16.433 39.34 16.633 ;
 RECT 39.116 16.433 39.172 16.633 ;
 RECT 38.276 16.433 38.332 16.633 ;
 RECT 38.108 16.433 38.164 16.633 ;
 RECT 38.612 16.433 38.668 16.633 ;
 RECT 38.444 16.433 38.5 16.633 ;
 RECT 37.604 16.433 37.66 16.633 ;
 RECT 37.436 16.433 37.492 16.633 ;
 RECT 37.94 16.433 37.996 16.633 ;
 RECT 37.772 16.433 37.828 16.633 ;
 RECT 36.932 16.433 36.988 16.633 ;
 RECT 36.764 16.433 36.82 16.633 ;
 RECT 37.268 16.433 37.324 16.633 ;
 RECT 37.1 16.433 37.156 16.633 ;
 RECT 36.26 16.433 36.316 16.633 ;
 RECT 36.092 16.433 36.148 16.633 ;
 RECT 36.596 16.433 36.652 16.633 ;
 RECT 36.428 16.433 36.484 16.633 ;
 RECT 35.588 16.433 35.644 16.633 ;
 RECT 35.42 16.433 35.476 16.633 ;
 RECT 35.252 16.433 35.308 16.633 ;
 RECT 35.924 16.433 35.98 16.633 ;
 RECT 35.756 16.433 35.812 16.633 ;
 RECT 40.124 17.2915 40.18 17.4915 ;
 RECT 39.62 17.2925 39.676 17.4925 ;
 RECT 39.452 17.2915 39.508 17.4915 ;
 RECT 39.956 17.106 40.012 17.306 ;
 RECT 39.788 17.2925 39.844 17.4925 ;
 RECT 38.948 17.2925 39.004 17.4925 ;
 RECT 38.78 17.2915 38.836 17.4915 ;
 RECT 39.284 17.106 39.34 17.306 ;
 RECT 39.116 17.2925 39.172 17.4925 ;
 RECT 38.276 17.2925 38.332 17.4925 ;
 RECT 38.108 17.2915 38.164 17.4915 ;
 RECT 38.612 17.106 38.668 17.306 ;
 RECT 38.444 17.2925 38.5 17.4925 ;
 RECT 37.604 17.2925 37.66 17.4925 ;
 RECT 37.436 17.2915 37.492 17.4915 ;
 RECT 37.94 17.106 37.996 17.306 ;
 RECT 37.772 17.2925 37.828 17.4925 ;
 RECT 36.932 17.2925 36.988 17.4925 ;
 RECT 36.764 17.2915 36.82 17.4915 ;
 RECT 37.268 17.106 37.324 17.306 ;
 RECT 37.1 17.2925 37.156 17.4925 ;
 RECT 36.26 17.2925 36.316 17.4925 ;
 RECT 36.092 17.2915 36.148 17.4915 ;
 RECT 36.596 17.106 36.652 17.306 ;
 RECT 36.428 17.2925 36.484 17.4925 ;
 RECT 35.588 17.2925 35.644 17.4925 ;
 RECT 35.42 17.2915 35.476 17.4915 ;
 RECT 35.252 17.106 35.308 17.306 ;
 RECT 35.924 17.106 35.98 17.306 ;
 RECT 35.756 17.2925 35.812 17.4925 ;
 END
 END vccdgt_1p0.gds1143
 PIN vccdgt_1p0.gds1144
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.162 15.679 45.202 15.879 ;
 END
 END vccdgt_1p0.gds1144
 PIN vccdgt_1p0.gds1145
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.49 15.679 44.53 15.879 ;
 END
 END vccdgt_1p0.gds1145
 PIN vccdgt_1p0.gds1146
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.818 15.679 43.858 15.879 ;
 END
 END vccdgt_1p0.gds1146
 PIN vccdgt_1p0.gds1147
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.146 15.679 43.186 15.879 ;
 END
 END vccdgt_1p0.gds1147
 PIN vccdgt_1p0.gds1148
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.474 15.679 42.514 15.879 ;
 END
 END vccdgt_1p0.gds1148
 PIN vccdgt_1p0.gds1149
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.802 15.679 41.842 15.879 ;
 END
 END vccdgt_1p0.gds1149
 PIN vccdgt_1p0.gds1150
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.13 15.679 41.17 15.879 ;
 END
 END vccdgt_1p0.gds1150
 PIN vccdgt_1p0.gds1151
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.742 17.5555 44.802 17.7555 ;
 END
 END vccdgt_1p0.gds1151
 PIN vccdgt_1p0.gds1152
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.07 17.5555 44.13 17.7555 ;
 END
 END vccdgt_1p0.gds1152
 PIN vccdgt_1p0.gds1153
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.398 17.5555 43.458 17.7555 ;
 END
 END vccdgt_1p0.gds1153
 PIN vccdgt_1p0.gds1154
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.726 17.5555 42.786 17.7555 ;
 END
 END vccdgt_1p0.gds1154
 PIN vccdgt_1p0.gds1155
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.054 17.5555 42.114 17.7555 ;
 END
 END vccdgt_1p0.gds1155
 PIN vccdgt_1p0.gds1156
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.382 17.5555 41.442 17.7555 ;
 END
 END vccdgt_1p0.gds1156
 PIN vccdgt_1p0.gds1157
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.29 17.5555 40.35 17.7555 ;
 END
 END vccdgt_1p0.gds1157
 PIN vccdgt_1p0.gds1158
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.982 18.16 41.022 18.36 ;
 END
 END vccdgt_1p0.gds1158
 PIN vccdgt_1p0.gds1159
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.71 17.915 40.75 18.115 ;
 END
 END vccdgt_1p0.gds1159
 PIN vccdgt_1p0.gds1160
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 45.164 18.127 45.22 18.327 ;
 RECT 44.66 18.127 44.716 18.327 ;
 RECT 44.492 18.127 44.548 18.327 ;
 RECT 44.828 18.127 44.884 18.327 ;
 RECT 44.996 18.127 45.052 18.327 ;
 RECT 43.988 18.127 44.044 18.327 ;
 RECT 43.82 18.127 43.876 18.327 ;
 RECT 44.156 18.127 44.212 18.327 ;
 RECT 44.324 18.127 44.38 18.327 ;
 RECT 43.316 18.127 43.372 18.327 ;
 RECT 43.148 18.127 43.204 18.327 ;
 RECT 43.484 18.127 43.54 18.327 ;
 RECT 43.652 18.127 43.708 18.327 ;
 RECT 42.644 18.127 42.7 18.327 ;
 RECT 42.476 18.127 42.532 18.327 ;
 RECT 42.812 18.127 42.868 18.327 ;
 RECT 42.98 18.127 43.036 18.327 ;
 RECT 41.972 18.127 42.028 18.327 ;
 RECT 41.804 18.127 41.86 18.327 ;
 RECT 42.14 18.127 42.196 18.327 ;
 RECT 42.308 18.127 42.364 18.327 ;
 RECT 41.3 18.127 41.356 18.327 ;
 RECT 41.132 18.127 41.188 18.327 ;
 RECT 41.468 18.127 41.524 18.327 ;
 RECT 41.636 18.127 41.692 18.327 ;
 RECT 40.544 18.127 40.6 18.327 ;
 RECT 40.376 18.127 40.432 18.327 ;
 RECT 44.744 16.433 44.8 16.633 ;
 RECT 44.576 16.433 44.632 16.633 ;
 RECT 45.08 16.433 45.136 16.633 ;
 RECT 44.912 16.433 44.968 16.633 ;
 RECT 44.072 16.433 44.128 16.633 ;
 RECT 43.904 16.433 43.96 16.633 ;
 RECT 44.408 16.433 44.464 16.633 ;
 RECT 44.24 16.433 44.296 16.633 ;
 RECT 43.4 16.433 43.456 16.633 ;
 RECT 43.232 16.433 43.288 16.633 ;
 RECT 43.736 16.433 43.792 16.633 ;
 RECT 43.568 16.433 43.624 16.633 ;
 RECT 42.728 16.433 42.784 16.633 ;
 RECT 42.56 16.433 42.616 16.633 ;
 RECT 43.064 16.433 43.12 16.633 ;
 RECT 42.896 16.433 42.952 16.633 ;
 RECT 42.056 16.433 42.112 16.633 ;
 RECT 41.888 16.433 41.944 16.633 ;
 RECT 42.392 16.433 42.448 16.633 ;
 RECT 42.224 16.433 42.28 16.633 ;
 RECT 41.384 16.433 41.44 16.633 ;
 RECT 41.216 16.433 41.272 16.633 ;
 RECT 41.048 16.433 41.104 16.633 ;
 RECT 41.72 16.433 41.776 16.633 ;
 RECT 41.552 16.433 41.608 16.633 ;
 RECT 40.628 16.433 40.684 16.633 ;
 RECT 40.46 16.433 40.516 16.633 ;
 RECT 40.292 16.433 40.348 16.633 ;
 RECT 40.88 16.434 40.936 16.634 ;
 RECT 44.744 17.2925 44.8 17.4925 ;
 RECT 44.576 17.2915 44.632 17.4915 ;
 RECT 45.08 17.106 45.136 17.306 ;
 RECT 44.912 17.2925 44.968 17.4925 ;
 RECT 44.072 17.2925 44.128 17.4925 ;
 RECT 43.904 17.2915 43.96 17.4915 ;
 RECT 44.408 17.106 44.464 17.306 ;
 RECT 44.24 17.2925 44.296 17.4925 ;
 RECT 43.4 17.2925 43.456 17.4925 ;
 RECT 43.232 17.2915 43.288 17.4915 ;
 RECT 43.736 17.106 43.792 17.306 ;
 RECT 43.568 17.2925 43.624 17.4925 ;
 RECT 42.728 17.2925 42.784 17.4925 ;
 RECT 42.56 17.2915 42.616 17.4915 ;
 RECT 43.064 17.106 43.12 17.306 ;
 RECT 42.896 17.2925 42.952 17.4925 ;
 RECT 42.056 17.2925 42.112 17.4925 ;
 RECT 41.888 17.2915 41.944 17.4915 ;
 RECT 42.392 17.106 42.448 17.306 ;
 RECT 42.224 17.2925 42.28 17.4925 ;
 RECT 41.384 17.2925 41.44 17.4925 ;
 RECT 41.216 17.2915 41.272 17.4915 ;
 RECT 41.048 17.106 41.104 17.306 ;
 RECT 41.72 17.106 41.776 17.306 ;
 RECT 41.552 17.2925 41.608 17.4925 ;
 RECT 40.628 17.106 40.684 17.306 ;
 RECT 40.46 17.2925 40.516 17.4925 ;
 RECT 40.292 17.2925 40.348 17.4925 ;
 RECT 40.964 17.2105 41.02 17.4105 ;
 RECT 40.712 17.3245 40.768 17.5245 ;
 END
 END vccdgt_1p0.gds1160
 PIN vccdgt_1p0.gds1161
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.866 15.447 47.922 15.647 ;
 END
 END vccdgt_1p0.gds1161
 PIN vccdgt_1p0.gds1162
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.834 15.679 45.874 15.879 ;
 END
 END vccdgt_1p0.gds1162
 PIN vccdgt_1p0.gds1163
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.446 18.348 47.502 18.548 ;
 END
 END vccdgt_1p0.gds1163
 PIN vccdgt_1p0.gds1164
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.97 18.185 50.03 18.385 ;
 END
 END vccdgt_1p0.gds1164
 PIN vccdgt_1p0.gds1165
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.626 17.2285 48.682 17.4285 ;
 END
 END vccdgt_1p0.gds1165
 PIN vccdgt_1p0.gds1166
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.29 18.664 49.33 18.864 ;
 END
 END vccdgt_1p0.gds1166
 PIN vccdgt_1p0.gds1167
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.086 17.5555 46.146 17.7555 ;
 END
 END vccdgt_1p0.gds1167
 PIN vccdgt_1p0.gds1168
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.414 17.5555 45.474 17.7555 ;
 END
 END vccdgt_1p0.gds1168
 PIN vccdgt_1p0.gds1169
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.418 18.5935 49.458 18.7935 ;
 END
 END vccdgt_1p0.gds1169
 PIN vccdgt_1p0.gds1170
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.606 18.5525 47.662 18.7525 ;
 END
 END vccdgt_1p0.gds1170
 PIN vccdgt_1p0.gds1171
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.266 18.266 47.342 18.466 ;
 END
 END vccdgt_1p0.gds1171
 PIN vccdgt_1p0.gds1172
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.106 18.154 48.182 18.354 ;
 END
 END vccdgt_1p0.gds1172
 PIN vccdgt_1p0.gds1173
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.87 17.3945 48.91 17.5945 ;
 END
 END vccdgt_1p0.gds1173
 PIN vccdgt_1p0.gds1174
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.286 18.2595 48.342 18.4595 ;
 END
 END vccdgt_1p0.gds1174
 PIN vccdgt_1p0.gds1175
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.062 18.084 49.102 18.284 ;
 END
 END vccdgt_1p0.gds1175
 PIN vccdgt_1p0.gds1176
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.626 17.757 49.686 17.957 ;
 END
 END vccdgt_1p0.gds1176
 PIN vccdgt_1p0.gds1177
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.782 18.3175 46.822 18.5175 ;
 END
 END vccdgt_1p0.gds1177
 PIN vccdgt_1p0.gds1178
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.134 17.965 50.18 18.165 ;
 END
 END vccdgt_1p0.gds1178
 PIN vccdgt_1p0.gds1179
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.506 18.4715 46.566 18.6715 ;
 END
 END vccdgt_1p0.gds1179
 PIN vccdgt_1p0.gds1180
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 46.004 18.127 46.06 18.327 ;
 RECT 45.836 18.127 45.892 18.327 ;
 RECT 46.172 18.127 46.228 18.327 ;
 RECT 46.34 18.127 46.396 18.327 ;
 RECT 45.332 18.127 45.388 18.327 ;
 RECT 45.5 18.127 45.556 18.327 ;
 RECT 45.668 18.127 45.724 18.327 ;
 RECT 47.768 16.434 47.824 16.634 ;
 RECT 46.928 16.434 46.984 16.634 ;
 RECT 47.6 16.434 47.656 16.634 ;
 RECT 47.264 16.434 47.32 16.634 ;
 RECT 47.096 16.434 47.152 16.634 ;
 RECT 48.272 16.434 48.328 16.634 ;
 RECT 48.104 16.434 48.16 16.634 ;
 RECT 49.28 16.434 49.336 16.634 ;
 RECT 49.112 16.434 49.168 16.634 ;
 RECT 48.944 16.434 49 16.634 ;
 RECT 48.776 16.431 48.832 16.631 ;
 RECT 48.608 16.434 48.664 16.634 ;
 RECT 50.204 16.434 50.26 16.634 ;
 RECT 49.868 16.434 49.924 16.634 ;
 RECT 49.7 16.434 49.756 16.634 ;
 RECT 49.532 16.434 49.588 16.634 ;
 RECT 46.088 16.433 46.144 16.633 ;
 RECT 45.92 16.433 45.976 16.633 ;
 RECT 46.424 16.433 46.48 16.633 ;
 RECT 46.256 16.433 46.312 16.633 ;
 RECT 45.416 16.433 45.472 16.633 ;
 RECT 45.248 16.433 45.304 16.633 ;
 RECT 45.752 16.433 45.808 16.633 ;
 RECT 45.584 16.433 45.64 16.633 ;
 RECT 47.768 17.63 47.824 17.83 ;
 RECT 46.928 17.63 46.984 17.83 ;
 RECT 48.44 17.742 48.496 17.942 ;
 RECT 46.592 17.3055 46.648 17.5055 ;
 RECT 46.76 17.533 46.816 17.733 ;
 RECT 48.272 17.6435 48.328 17.8435 ;
 RECT 48.104 17.5755 48.16 17.7755 ;
 RECT 47.936 17.472 47.992 17.672 ;
 RECT 50.204 19.157 50.26 19.357 ;
 RECT 48.104 19.04 48.16 19.24 ;
 RECT 48.86 19.157 48.916 19.357 ;
 RECT 46.508 16.183 46.564 16.383 ;
 RECT 47.432 16.63 47.488 16.83 ;
 RECT 48.86 20.417 48.916 20.617 ;
 RECT 49.028 19.984 49.084 20.184 ;
 RECT 49.868 20.06 49.924 20.26 ;
 RECT 48.104 20.3 48.16 20.5 ;
 RECT 49.616 20.312 49.672 20.512 ;
 RECT 49.364 20.399 49.42 20.599 ;
 RECT 48.692 20.417 48.748 20.617 ;
 RECT 50.204 20.417 50.26 20.617 ;
 RECT 48.524 20.404 48.58 20.604 ;
 RECT 49.028 18.724 49.084 18.924 ;
 RECT 49.868 18.8 49.924 19 ;
 RECT 49.616 19.052 49.672 19.252 ;
 RECT 50.036 19.22 50.092 19.42 ;
 RECT 48.944 17.533 49 17.733 ;
 RECT 48.608 17.5895 48.664 17.7895 ;
 RECT 48.776 17.6715 48.832 17.8715 ;
 RECT 49.112 17.533 49.168 17.733 ;
 RECT 49.28 17.5895 49.336 17.7895 ;
 RECT 49.784 17.6715 49.84 17.8715 ;
 RECT 49.448 17.601 49.504 17.801 ;
 RECT 49.616 17.5895 49.672 17.7895 ;
 RECT 50.12 17.533 50.176 17.733 ;
 RECT 49.952 17.533 50.008 17.733 ;
 RECT 49.364 19.139 49.42 19.339 ;
 RECT 48.692 19.157 48.748 19.357 ;
 RECT 48.524 19.144 48.58 19.344 ;
 RECT 46.088 17.2925 46.144 17.4925 ;
 RECT 45.92 17.2915 45.976 17.4915 ;
 RECT 46.424 17.106 46.48 17.306 ;
 RECT 46.256 17.2925 46.312 17.4925 ;
 RECT 45.416 17.2925 45.472 17.4925 ;
 RECT 45.248 17.2915 45.304 17.4915 ;
 RECT 45.752 17.106 45.808 17.306 ;
 RECT 45.584 17.2925 45.64 17.4925 ;
 END
 END vccdgt_1p0.gds1180
 PIN vccdgt_1p0.gds1181
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.074 15.679 55.114 15.879 ;
 END
 END vccdgt_1p0.gds1181
 PIN vccdgt_1p0.gds1182
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.402 15.679 54.442 15.879 ;
 END
 END vccdgt_1p0.gds1182
 PIN vccdgt_1p0.gds1183
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.73 15.679 53.77 15.879 ;
 END
 END vccdgt_1p0.gds1183
 PIN vccdgt_1p0.gds1184
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.058 15.679 53.098 15.879 ;
 END
 END vccdgt_1p0.gds1184
 PIN vccdgt_1p0.gds1185
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.386 15.679 52.426 15.879 ;
 END
 END vccdgt_1p0.gds1185
 PIN vccdgt_1p0.gds1186
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 19.666 50.674 19.866 ;
 END
 END vccdgt_1p0.gds1186
 PIN vccdgt_1p0.gds1187
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.942 19.5775 50.998 19.7775 ;
 END
 END vccdgt_1p0.gds1187
 PIN vccdgt_1p0.gds1188
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.778 18.911 50.838 19.111 ;
 END
 END vccdgt_1p0.gds1188
 PIN vccdgt_1p0.gds1189
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.122 19.3865 51.178 19.5865 ;
 END
 END vccdgt_1p0.gds1189
 PIN vccdgt_1p0.gds1190
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.654 17.5555 54.714 17.7555 ;
 END
 END vccdgt_1p0.gds1190
 PIN vccdgt_1p0.gds1191
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.982 17.5555 54.042 17.7555 ;
 END
 END vccdgt_1p0.gds1191
 PIN vccdgt_1p0.gds1192
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.31 17.5555 53.37 17.7555 ;
 END
 END vccdgt_1p0.gds1192
 PIN vccdgt_1p0.gds1193
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.638 17.5555 52.698 17.7555 ;
 END
 END vccdgt_1p0.gds1193
 PIN vccdgt_1p0.gds1194
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.442 18.1605 51.518 18.3605 ;
 END
 END vccdgt_1p0.gds1194
 PIN vccdgt_1p0.gds1195
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 17.697 50.674 17.897 ;
 END
 END vccdgt_1p0.gds1195
 PIN vccdgt_1p0.gds1196
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.218 18.2535 52.278 18.4535 ;
 END
 END vccdgt_1p0.gds1196
 PIN vccdgt_1p0.gds1197
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.962 19.4835 52.002 19.6835 ;
 END
 END vccdgt_1p0.gds1197
 PIN vccdgt_1p0.gds1198
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.282 17.8845 51.338 18.0845 ;
 END
 END vccdgt_1p0.gds1198
 PIN vccdgt_1p0.gds1199
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.702 17.845 51.758 18.045 ;
 END
 END vccdgt_1p0.gds1199
 PIN vccdgt_1p0.gds1200
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 55.076 18.127 55.132 18.327 ;
 RECT 54.572 18.127 54.628 18.327 ;
 RECT 54.404 18.127 54.46 18.327 ;
 RECT 54.74 18.127 54.796 18.327 ;
 RECT 54.908 18.127 54.964 18.327 ;
 RECT 53.9 18.127 53.956 18.327 ;
 RECT 53.732 18.127 53.788 18.327 ;
 RECT 54.068 18.127 54.124 18.327 ;
 RECT 54.236 18.127 54.292 18.327 ;
 RECT 53.228 18.127 53.284 18.327 ;
 RECT 53.06 18.127 53.116 18.327 ;
 RECT 53.396 18.127 53.452 18.327 ;
 RECT 53.564 18.127 53.62 18.327 ;
 RECT 52.556 18.127 52.612 18.327 ;
 RECT 52.388 18.127 52.444 18.327 ;
 RECT 52.892 18.127 52.948 18.327 ;
 RECT 52.724 18.127 52.78 18.327 ;
 RECT 55.16 16.433 55.216 16.633 ;
 RECT 54.656 16.433 54.712 16.633 ;
 RECT 54.488 16.433 54.544 16.633 ;
 RECT 54.992 16.433 55.048 16.633 ;
 RECT 54.824 16.433 54.88 16.633 ;
 RECT 53.984 16.433 54.04 16.633 ;
 RECT 53.816 16.433 53.872 16.633 ;
 RECT 54.32 16.433 54.376 16.633 ;
 RECT 54.152 16.433 54.208 16.633 ;
 RECT 50.876 16.434 50.932 16.634 ;
 RECT 50.708 16.434 50.764 16.634 ;
 RECT 50.54 16.434 50.596 16.634 ;
 RECT 50.372 16.434 50.428 16.634 ;
 RECT 51.38 16.471 51.436 16.653 ;
 RECT 51.128 16.471 51.184 16.653 ;
 RECT 51.716 16.435 51.772 16.635 ;
 RECT 53.312 16.433 53.368 16.633 ;
 RECT 53.144 16.433 53.2 16.633 ;
 RECT 53.648 16.433 53.704 16.633 ;
 RECT 53.48 16.433 53.536 16.633 ;
 RECT 52.64 16.433 52.696 16.633 ;
 RECT 52.472 16.433 52.528 16.633 ;
 RECT 52.304 16.433 52.36 16.633 ;
 RECT 52.976 16.433 53.032 16.633 ;
 RECT 52.808 16.433 52.864 16.633 ;
 RECT 52.136 17.783 52.192 17.983 ;
 RECT 52.22 15.621 52.276 15.821 ;
 RECT 55.16 17.2915 55.216 17.4915 ;
 RECT 54.656 17.2925 54.712 17.4925 ;
 RECT 54.488 17.2915 54.544 17.4915 ;
 RECT 54.992 17.106 55.048 17.306 ;
 RECT 54.824 17.2925 54.88 17.4925 ;
 RECT 53.984 17.2925 54.04 17.4925 ;
 RECT 53.816 17.2915 53.872 17.4915 ;
 RECT 54.32 17.106 54.376 17.306 ;
 RECT 54.152 17.2925 54.208 17.4925 ;
 RECT 50.96 17.533 51.016 17.733 ;
 RECT 50.792 17.533 50.848 17.733 ;
 RECT 50.624 17.533 50.68 17.733 ;
 RECT 50.456 17.533 50.512 17.733 ;
 RECT 50.288 17.533 50.344 17.733 ;
 RECT 51.8 17.4855 51.856 17.6855 ;
 RECT 51.464 17.5645 51.52 17.7645 ;
 RECT 51.128 17.498 51.184 17.698 ;
 RECT 51.632 17.5645 51.688 17.7645 ;
 RECT 51.296 17.4855 51.352 17.6855 ;
 RECT 51.968 17.4855 52.024 17.6855 ;
 RECT 53.312 17.2925 53.368 17.4925 ;
 RECT 53.144 17.2915 53.2 17.4915 ;
 RECT 53.648 17.106 53.704 17.306 ;
 RECT 53.48 17.2925 53.536 17.4925 ;
 RECT 52.64 17.2925 52.696 17.4925 ;
 RECT 52.472 17.2915 52.528 17.4915 ;
 RECT 52.304 17.106 52.36 17.306 ;
 RECT 52.976 17.106 53.032 17.306 ;
 RECT 52.808 17.2925 52.864 17.4925 ;
 END
 END vccdgt_1p0.gds1200
 PIN vccdgt_1p0.gds1201
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.182 15.679 58.222 15.879 ;
 END
 END vccdgt_1p0.gds1201
 PIN vccdgt_1p0.gds1202
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.09 15.679 57.13 15.879 ;
 END
 END vccdgt_1p0.gds1202
 PIN vccdgt_1p0.gds1203
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.198 15.679 60.238 15.879 ;
 END
 END vccdgt_1p0.gds1203
 PIN vccdgt_1p0.gds1204
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.526 15.679 59.566 15.879 ;
 END
 END vccdgt_1p0.gds1204
 PIN vccdgt_1p0.gds1205
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.854 15.679 58.894 15.879 ;
 END
 END vccdgt_1p0.gds1205
 PIN vccdgt_1p0.gds1206
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.418 15.679 56.458 15.879 ;
 END
 END vccdgt_1p0.gds1206
 PIN vccdgt_1p0.gds1207
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.746 15.679 55.786 15.879 ;
 END
 END vccdgt_1p0.gds1207
 PIN vccdgt_1p0.gds1208
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.778 17.5555 59.838 17.7555 ;
 END
 END vccdgt_1p0.gds1208
 PIN vccdgt_1p0.gds1209
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.106 17.5555 59.166 17.7555 ;
 END
 END vccdgt_1p0.gds1209
 PIN vccdgt_1p0.gds1210
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.434 17.5555 58.494 17.7555 ;
 END
 END vccdgt_1p0.gds1210
 PIN vccdgt_1p0.gds1211
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.342 17.5555 57.402 17.7555 ;
 END
 END vccdgt_1p0.gds1211
 PIN vccdgt_1p0.gds1212
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.67 17.5555 56.73 17.7555 ;
 END
 END vccdgt_1p0.gds1212
 PIN vccdgt_1p0.gds1213
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.998 17.5555 56.058 17.7555 ;
 END
 END vccdgt_1p0.gds1213
 PIN vccdgt_1p0.gds1214
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.326 17.5555 55.386 17.7555 ;
 END
 END vccdgt_1p0.gds1214
 PIN vccdgt_1p0.gds1215
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.034 18.16 58.074 18.36 ;
 END
 END vccdgt_1p0.gds1215
 PIN vccdgt_1p0.gds1216
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.762 17.915 57.802 18.115 ;
 END
 END vccdgt_1p0.gds1216
 PIN vccdgt_1p0.gds1217
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 60.2 18.127 60.256 18.327 ;
 RECT 59.696 18.127 59.752 18.327 ;
 RECT 59.528 18.127 59.584 18.327 ;
 RECT 59.864 18.127 59.92 18.327 ;
 RECT 60.032 18.127 60.088 18.327 ;
 RECT 59.024 18.127 59.08 18.327 ;
 RECT 58.856 18.127 58.912 18.327 ;
 RECT 59.192 18.127 59.248 18.327 ;
 RECT 59.36 18.127 59.416 18.327 ;
 RECT 58.352 18.127 58.408 18.327 ;
 RECT 58.184 18.127 58.24 18.327 ;
 RECT 58.52 18.127 58.576 18.327 ;
 RECT 58.688 18.127 58.744 18.327 ;
 RECT 57.26 18.127 57.316 18.327 ;
 RECT 57.092 18.127 57.148 18.327 ;
 RECT 57.428 18.127 57.484 18.327 ;
 RECT 57.596 18.127 57.652 18.327 ;
 RECT 56.588 18.127 56.644 18.327 ;
 RECT 56.42 18.127 56.476 18.327 ;
 RECT 56.756 18.127 56.812 18.327 ;
 RECT 56.924 18.127 56.98 18.327 ;
 RECT 55.916 18.127 55.972 18.327 ;
 RECT 55.748 18.127 55.804 18.327 ;
 RECT 56.084 18.127 56.14 18.327 ;
 RECT 56.252 18.127 56.308 18.327 ;
 RECT 55.244 18.127 55.3 18.327 ;
 RECT 55.412 18.127 55.468 18.327 ;
 RECT 55.58 18.127 55.636 18.327 ;
 RECT 59.78 16.433 59.836 16.633 ;
 RECT 59.612 16.433 59.668 16.633 ;
 RECT 60.116 16.433 60.172 16.633 ;
 RECT 59.948 16.433 60.004 16.633 ;
 RECT 59.108 16.433 59.164 16.633 ;
 RECT 58.94 16.433 58.996 16.633 ;
 RECT 59.444 16.433 59.5 16.633 ;
 RECT 59.276 16.433 59.332 16.633 ;
 RECT 58.436 16.433 58.492 16.633 ;
 RECT 58.268 16.433 58.324 16.633 ;
 RECT 58.1 16.433 58.156 16.633 ;
 RECT 58.772 16.433 58.828 16.633 ;
 RECT 58.604 16.433 58.66 16.633 ;
 RECT 57.344 16.433 57.4 16.633 ;
 RECT 57.176 16.433 57.232 16.633 ;
 RECT 57.68 16.433 57.736 16.633 ;
 RECT 57.512 16.433 57.568 16.633 ;
 RECT 56.672 16.433 56.728 16.633 ;
 RECT 56.504 16.433 56.56 16.633 ;
 RECT 57.008 16.433 57.064 16.633 ;
 RECT 56.84 16.433 56.896 16.633 ;
 RECT 56 16.433 56.056 16.633 ;
 RECT 55.832 16.433 55.888 16.633 ;
 RECT 56.336 16.433 56.392 16.633 ;
 RECT 56.168 16.433 56.224 16.633 ;
 RECT 55.328 16.433 55.384 16.633 ;
 RECT 55.664 16.433 55.72 16.633 ;
 RECT 55.496 16.433 55.552 16.633 ;
 RECT 57.932 16.434 57.988 16.634 ;
 RECT 58.016 17.2105 58.072 17.4105 ;
 RECT 57.764 17.3245 57.82 17.5245 ;
 RECT 59.78 17.2925 59.836 17.4925 ;
 RECT 59.612 17.2915 59.668 17.4915 ;
 RECT 60.116 17.106 60.172 17.306 ;
 RECT 59.948 17.2925 60.004 17.4925 ;
 RECT 59.108 17.2925 59.164 17.4925 ;
 RECT 58.94 17.2915 58.996 17.4915 ;
 RECT 59.444 17.106 59.5 17.306 ;
 RECT 59.276 17.2925 59.332 17.4925 ;
 RECT 58.436 17.2925 58.492 17.4925 ;
 RECT 58.268 17.2915 58.324 17.4915 ;
 RECT 58.1 17.106 58.156 17.306 ;
 RECT 58.772 17.106 58.828 17.306 ;
 RECT 58.604 17.2925 58.66 17.4925 ;
 RECT 57.344 17.2925 57.4 17.4925 ;
 RECT 57.176 17.2915 57.232 17.4915 ;
 RECT 57.68 17.106 57.736 17.306 ;
 RECT 57.512 17.2925 57.568 17.4925 ;
 RECT 56.672 17.2925 56.728 17.4925 ;
 RECT 56.504 17.2915 56.56 17.4915 ;
 RECT 57.008 17.106 57.064 17.306 ;
 RECT 56.84 17.2925 56.896 17.4925 ;
 RECT 56 17.2925 56.056 17.4925 ;
 RECT 55.832 17.2915 55.888 17.4915 ;
 RECT 56.336 17.106 56.392 17.306 ;
 RECT 56.168 17.2925 56.224 17.4925 ;
 RECT 55.328 17.2925 55.384 17.4925 ;
 RECT 55.664 17.106 55.72 17.306 ;
 RECT 55.496 17.2925 55.552 17.4925 ;
 END
 END vccdgt_1p0.gds1217
 PIN vccdgt_1p0.gds1218
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.918 15.447 64.974 15.647 ;
 END
 END vccdgt_1p0.gds1218
 PIN vccdgt_1p0.gds1219
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.886 15.679 62.926 15.879 ;
 END
 END vccdgt_1p0.gds1219
 PIN vccdgt_1p0.gds1220
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.214 15.679 62.254 15.879 ;
 END
 END vccdgt_1p0.gds1220
 PIN vccdgt_1p0.gds1221
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.542 15.679 61.582 15.879 ;
 END
 END vccdgt_1p0.gds1221
 PIN vccdgt_1p0.gds1222
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.87 15.679 60.91 15.879 ;
 END
 END vccdgt_1p0.gds1222
 PIN vccdgt_1p0.gds1223
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.498 18.348 64.554 18.548 ;
 END
 END vccdgt_1p0.gds1223
 PIN vccdgt_1p0.gds1224
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.138 17.5555 63.198 17.7555 ;
 END
 END vccdgt_1p0.gds1224
 PIN vccdgt_1p0.gds1225
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.466 17.5555 62.526 17.7555 ;
 END
 END vccdgt_1p0.gds1225
 PIN vccdgt_1p0.gds1226
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.794 17.5555 61.854 17.7555 ;
 END
 END vccdgt_1p0.gds1226
 PIN vccdgt_1p0.gds1227
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.122 17.5555 61.182 17.7555 ;
 END
 END vccdgt_1p0.gds1227
 PIN vccdgt_1p0.gds1228
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.45 17.5555 60.51 17.7555 ;
 END
 END vccdgt_1p0.gds1228
 PIN vccdgt_1p0.gds1229
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.658 18.5525 64.714 18.7525 ;
 END
 END vccdgt_1p0.gds1229
 PIN vccdgt_1p0.gds1230
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.318 18.266 64.394 18.466 ;
 END
 END vccdgt_1p0.gds1230
 PIN vccdgt_1p0.gds1231
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.834 18.3175 63.874 18.5175 ;
 END
 END vccdgt_1p0.gds1231
 PIN vccdgt_1p0.gds1232
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.158 18.154 65.234 18.354 ;
 END
 END vccdgt_1p0.gds1232
 PIN vccdgt_1p0.gds1233
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.558 18.4715 63.618 18.6715 ;
 END
 END vccdgt_1p0.gds1233
 PIN vccdgt_1p0.gds1234
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 63.056 18.127 63.112 18.327 ;
 RECT 62.888 18.127 62.944 18.327 ;
 RECT 63.224 18.127 63.28 18.327 ;
 RECT 63.392 18.127 63.448 18.327 ;
 RECT 62.384 18.127 62.44 18.327 ;
 RECT 62.216 18.127 62.272 18.327 ;
 RECT 62.552 18.127 62.608 18.327 ;
 RECT 62.72 18.127 62.776 18.327 ;
 RECT 61.712 18.127 61.768 18.327 ;
 RECT 61.544 18.127 61.6 18.327 ;
 RECT 61.88 18.127 61.936 18.327 ;
 RECT 62.048 18.127 62.104 18.327 ;
 RECT 61.04 18.127 61.096 18.327 ;
 RECT 60.872 18.127 60.928 18.327 ;
 RECT 61.208 18.127 61.264 18.327 ;
 RECT 61.376 18.127 61.432 18.327 ;
 RECT 60.536 18.127 60.592 18.327 ;
 RECT 60.704 18.127 60.76 18.327 ;
 RECT 60.368 18.127 60.424 18.327 ;
 RECT 64.82 16.434 64.876 16.634 ;
 RECT 63.98 16.434 64.036 16.634 ;
 RECT 64.652 16.434 64.708 16.634 ;
 RECT 64.316 16.434 64.372 16.634 ;
 RECT 64.148 16.434 64.204 16.634 ;
 RECT 65.156 16.434 65.212 16.634 ;
 RECT 63.14 16.433 63.196 16.633 ;
 RECT 62.972 16.433 63.028 16.633 ;
 RECT 63.476 16.433 63.532 16.633 ;
 RECT 63.308 16.433 63.364 16.633 ;
 RECT 62.468 16.433 62.524 16.633 ;
 RECT 62.3 16.433 62.356 16.633 ;
 RECT 62.804 16.433 62.86 16.633 ;
 RECT 62.636 16.433 62.692 16.633 ;
 RECT 61.796 16.433 61.852 16.633 ;
 RECT 61.628 16.433 61.684 16.633 ;
 RECT 62.132 16.433 62.188 16.633 ;
 RECT 61.964 16.433 62.02 16.633 ;
 RECT 61.124 16.433 61.18 16.633 ;
 RECT 60.956 16.433 61.012 16.633 ;
 RECT 61.46 16.433 61.516 16.633 ;
 RECT 61.292 16.433 61.348 16.633 ;
 RECT 60.452 16.433 60.508 16.633 ;
 RECT 60.788 16.433 60.844 16.633 ;
 RECT 60.62 16.433 60.676 16.633 ;
 RECT 60.284 16.433 60.34 16.633 ;
 RECT 64.82 17.63 64.876 17.83 ;
 RECT 63.98 17.63 64.036 17.83 ;
 RECT 63.644 17.3055 63.7 17.5055 ;
 RECT 63.812 17.533 63.868 17.733 ;
 RECT 65.156 17.5755 65.212 17.7755 ;
 RECT 64.988 17.472 65.044 17.672 ;
 RECT 65.156 20.3 65.212 20.5 ;
 RECT 65.156 19.04 65.212 19.24 ;
 RECT 63.56 16.183 63.616 16.383 ;
 RECT 64.484 16.63 64.54 16.83 ;
 RECT 63.14 17.2925 63.196 17.4925 ;
 RECT 62.972 17.2915 63.028 17.4915 ;
 RECT 63.476 17.106 63.532 17.306 ;
 RECT 63.308 17.2925 63.364 17.4925 ;
 RECT 62.468 17.2925 62.524 17.4925 ;
 RECT 62.3 17.2915 62.356 17.4915 ;
 RECT 62.804 17.106 62.86 17.306 ;
 RECT 62.636 17.2925 62.692 17.4925 ;
 RECT 61.796 17.2925 61.852 17.4925 ;
 RECT 61.628 17.2915 61.684 17.4915 ;
 RECT 62.132 17.106 62.188 17.306 ;
 RECT 61.964 17.2925 62.02 17.4925 ;
 RECT 61.124 17.2925 61.18 17.4925 ;
 RECT 60.956 17.2915 61.012 17.4915 ;
 RECT 61.46 17.106 61.516 17.306 ;
 RECT 61.292 17.2925 61.348 17.4925 ;
 RECT 60.452 17.2925 60.508 17.4925 ;
 RECT 60.788 17.106 60.844 17.306 ;
 RECT 60.62 17.2925 60.676 17.4925 ;
 RECT 60.284 17.2915 60.34 17.4915 ;
 END
 END vccdgt_1p0.gds1234
 PIN vccdgt_1p0.gds1235
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 19.666 67.726 19.866 ;
 END
 END vccdgt_1p0.gds1235
 PIN vccdgt_1p0.gds1236
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.678 17.2285 65.734 17.4285 ;
 END
 END vccdgt_1p0.gds1236
 PIN vccdgt_1p0.gds1237
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.022 18.185 67.082 18.385 ;
 END
 END vccdgt_1p0.gds1237
 PIN vccdgt_1p0.gds1238
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.342 18.664 66.382 18.864 ;
 END
 END vccdgt_1p0.gds1238
 PIN vccdgt_1p0.gds1239
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.11 15.679 70.15 15.879 ;
 END
 END vccdgt_1p0.gds1239
 PIN vccdgt_1p0.gds1240
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.438 15.679 69.478 15.879 ;
 END
 END vccdgt_1p0.gds1240
 PIN vccdgt_1p0.gds1241
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.994 19.5775 68.05 19.7775 ;
 END
 END vccdgt_1p0.gds1241
 PIN vccdgt_1p0.gds1242
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.83 18.911 67.89 19.111 ;
 END
 END vccdgt_1p0.gds1242
 PIN vccdgt_1p0.gds1243
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.174 19.3865 68.23 19.5865 ;
 END
 END vccdgt_1p0.gds1243
 PIN vccdgt_1p0.gds1244
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.69 17.5555 69.75 17.7555 ;
 END
 END vccdgt_1p0.gds1244
 PIN vccdgt_1p0.gds1245
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.494 18.1605 68.57 18.3605 ;
 END
 END vccdgt_1p0.gds1245
 PIN vccdgt_1p0.gds1246
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.47 18.5935 66.51 18.7935 ;
 END
 END vccdgt_1p0.gds1246
 PIN vccdgt_1p0.gds1247
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.922 17.3945 65.962 17.5945 ;
 END
 END vccdgt_1p0.gds1247
 PIN vccdgt_1p0.gds1248
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.338 18.2595 65.394 18.4595 ;
 END
 END vccdgt_1p0.gds1248
 PIN vccdgt_1p0.gds1249
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.27 18.2535 69.33 18.4535 ;
 END
 END vccdgt_1p0.gds1249
 PIN vccdgt_1p0.gds1250
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.014 19.4835 69.054 19.6835 ;
 END
 END vccdgt_1p0.gds1250
 PIN vccdgt_1p0.gds1251
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.334 17.8845 68.39 18.0845 ;
 END
 END vccdgt_1p0.gds1251
 PIN vccdgt_1p0.gds1252
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.114 18.084 66.154 18.284 ;
 END
 END vccdgt_1p0.gds1252
 PIN vccdgt_1p0.gds1253
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.754 17.845 68.81 18.045 ;
 END
 END vccdgt_1p0.gds1253
 PIN vccdgt_1p0.gds1254
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.678 17.757 66.738 17.957 ;
 END
 END vccdgt_1p0.gds1254
 PIN vccdgt_1p0.gds1255
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 17.697 67.726 17.897 ;
 END
 END vccdgt_1p0.gds1255
 PIN vccdgt_1p0.gds1256
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.186 17.965 67.232 18.165 ;
 END
 END vccdgt_1p0.gds1256
 PIN vccdgt_1p0.gds1257
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 70.112 18.127 70.168 18.327 ;
 RECT 69.608 18.127 69.664 18.327 ;
 RECT 69.44 18.127 69.496 18.327 ;
 RECT 69.944 18.127 70 18.327 ;
 RECT 69.776 18.127 69.832 18.327 ;
 RECT 65.324 16.434 65.38 16.634 ;
 RECT 66.332 16.434 66.388 16.634 ;
 RECT 66.164 16.434 66.22 16.634 ;
 RECT 65.996 16.434 66.052 16.634 ;
 RECT 65.828 16.431 65.884 16.631 ;
 RECT 65.66 16.434 65.716 16.634 ;
 RECT 67.256 16.434 67.312 16.634 ;
 RECT 66.92 16.434 66.976 16.634 ;
 RECT 66.752 16.434 66.808 16.634 ;
 RECT 66.584 16.434 66.64 16.634 ;
 RECT 67.928 16.434 67.984 16.634 ;
 RECT 67.76 16.434 67.816 16.634 ;
 RECT 67.592 16.434 67.648 16.634 ;
 RECT 67.424 16.434 67.48 16.634 ;
 RECT 68.432 16.471 68.488 16.653 ;
 RECT 68.18 16.471 68.236 16.653 ;
 RECT 68.768 16.435 68.824 16.635 ;
 RECT 70.196 16.433 70.252 16.633 ;
 RECT 69.692 16.433 69.748 16.633 ;
 RECT 69.524 16.433 69.58 16.633 ;
 RECT 69.356 16.433 69.412 16.633 ;
 RECT 70.028 16.433 70.084 16.633 ;
 RECT 69.86 16.433 69.916 16.633 ;
 RECT 65.492 17.742 65.548 17.942 ;
 RECT 69.188 17.783 69.244 17.983 ;
 RECT 65.324 17.6435 65.38 17.8435 ;
 RECT 67.256 19.157 67.312 19.357 ;
 RECT 65.912 19.157 65.968 19.357 ;
 RECT 65.912 20.417 65.968 20.617 ;
 RECT 66.08 19.984 66.136 20.184 ;
 RECT 66.92 20.06 66.976 20.26 ;
 RECT 66.668 20.312 66.724 20.512 ;
 RECT 66.416 20.399 66.472 20.599 ;
 RECT 65.744 20.417 65.8 20.617 ;
 RECT 67.256 20.417 67.312 20.617 ;
 RECT 65.576 20.404 65.632 20.604 ;
 RECT 66.08 18.724 66.136 18.924 ;
 RECT 66.92 18.8 66.976 19 ;
 RECT 66.668 19.052 66.724 19.252 ;
 RECT 67.088 19.22 67.144 19.42 ;
 RECT 66.416 19.139 66.472 19.339 ;
 RECT 65.744 19.157 65.8 19.357 ;
 RECT 65.576 19.144 65.632 19.344 ;
 RECT 69.272 15.621 69.328 15.821 ;
 RECT 65.996 17.533 66.052 17.733 ;
 RECT 65.66 17.5895 65.716 17.7895 ;
 RECT 65.828 17.6715 65.884 17.8715 ;
 RECT 66.164 17.533 66.22 17.733 ;
 RECT 66.332 17.5895 66.388 17.7895 ;
 RECT 68.012 17.533 68.068 17.733 ;
 RECT 66.836 17.6715 66.892 17.8715 ;
 RECT 66.5 17.601 66.556 17.801 ;
 RECT 66.668 17.5895 66.724 17.7895 ;
 RECT 67.172 17.533 67.228 17.733 ;
 RECT 67.004 17.533 67.06 17.733 ;
 RECT 67.844 17.533 67.9 17.733 ;
 RECT 67.676 17.533 67.732 17.733 ;
 RECT 67.508 17.533 67.564 17.733 ;
 RECT 67.34 17.533 67.396 17.733 ;
 RECT 68.852 17.4855 68.908 17.6855 ;
 RECT 68.516 17.5645 68.572 17.7645 ;
 RECT 68.18 17.498 68.236 17.698 ;
 RECT 68.684 17.5645 68.74 17.7645 ;
 RECT 68.348 17.4855 68.404 17.6855 ;
 RECT 69.02 17.4855 69.076 17.6855 ;
 RECT 70.196 17.2915 70.252 17.4915 ;
 RECT 69.692 17.2925 69.748 17.4925 ;
 RECT 69.524 17.2915 69.58 17.4915 ;
 RECT 69.356 17.106 69.412 17.306 ;
 RECT 70.028 17.106 70.084 17.306 ;
 RECT 69.86 17.2925 69.916 17.4925 ;
 END
 END vccdgt_1p0.gds1257
 PIN vccdgt_1p0.gds1258
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.142 15.679 74.182 15.879 ;
 END
 END vccdgt_1p0.gds1258
 PIN vccdgt_1p0.gds1259
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.47 15.679 73.51 15.879 ;
 END
 END vccdgt_1p0.gds1259
 PIN vccdgt_1p0.gds1260
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.798 15.679 72.838 15.879 ;
 END
 END vccdgt_1p0.gds1260
 PIN vccdgt_1p0.gds1261
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.126 15.679 72.166 15.879 ;
 END
 END vccdgt_1p0.gds1261
 PIN vccdgt_1p0.gds1262
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.454 15.679 71.494 15.879 ;
 END
 END vccdgt_1p0.gds1262
 PIN vccdgt_1p0.gds1263
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.782 15.679 70.822 15.879 ;
 END
 END vccdgt_1p0.gds1263
 PIN vccdgt_1p0.gds1264
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.394 17.5555 74.454 17.7555 ;
 END
 END vccdgt_1p0.gds1264
 PIN vccdgt_1p0.gds1265
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.722 17.5555 73.782 17.7555 ;
 END
 END vccdgt_1p0.gds1265
 PIN vccdgt_1p0.gds1266
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.05 17.5555 73.11 17.7555 ;
 END
 END vccdgt_1p0.gds1266
 PIN vccdgt_1p0.gds1267
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.378 17.5555 72.438 17.7555 ;
 END
 END vccdgt_1p0.gds1267
 PIN vccdgt_1p0.gds1268
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.706 17.5555 71.766 17.7555 ;
 END
 END vccdgt_1p0.gds1268
 PIN vccdgt_1p0.gds1269
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.034 17.5555 71.094 17.7555 ;
 END
 END vccdgt_1p0.gds1269
 PIN vccdgt_1p0.gds1270
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.362 17.5555 70.422 17.7555 ;
 END
 END vccdgt_1p0.gds1270
 PIN vccdgt_1p0.gds1271
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 74.312 18.127 74.368 18.327 ;
 RECT 74.144 18.127 74.2 18.327 ;
 RECT 74.48 18.127 74.536 18.327 ;
 RECT 74.648 18.127 74.704 18.327 ;
 RECT 73.64 18.127 73.696 18.327 ;
 RECT 73.472 18.127 73.528 18.327 ;
 RECT 73.808 18.127 73.864 18.327 ;
 RECT 73.976 18.127 74.032 18.327 ;
 RECT 72.968 18.127 73.024 18.327 ;
 RECT 72.8 18.127 72.856 18.327 ;
 RECT 73.136 18.127 73.192 18.327 ;
 RECT 73.304 18.127 73.36 18.327 ;
 RECT 72.296 18.127 72.352 18.327 ;
 RECT 72.128 18.127 72.184 18.327 ;
 RECT 72.464 18.127 72.52 18.327 ;
 RECT 72.632 18.127 72.688 18.327 ;
 RECT 71.624 18.127 71.68 18.327 ;
 RECT 71.456 18.127 71.512 18.327 ;
 RECT 71.792 18.127 71.848 18.327 ;
 RECT 71.96 18.127 72.016 18.327 ;
 RECT 70.952 18.127 71.008 18.327 ;
 RECT 70.784 18.127 70.84 18.327 ;
 RECT 71.12 18.127 71.176 18.327 ;
 RECT 71.288 18.127 71.344 18.327 ;
 RECT 70.28 18.127 70.336 18.327 ;
 RECT 70.448 18.127 70.504 18.327 ;
 RECT 70.616 18.127 70.672 18.327 ;
 RECT 74.396 16.433 74.452 16.633 ;
 RECT 74.228 16.433 74.284 16.633 ;
 RECT 74.732 16.433 74.788 16.633 ;
 RECT 74.564 16.433 74.62 16.633 ;
 RECT 73.724 16.433 73.78 16.633 ;
 RECT 73.556 16.433 73.612 16.633 ;
 RECT 74.06 16.433 74.116 16.633 ;
 RECT 73.892 16.433 73.948 16.633 ;
 RECT 73.052 16.433 73.108 16.633 ;
 RECT 72.884 16.433 72.94 16.633 ;
 RECT 73.388 16.433 73.444 16.633 ;
 RECT 73.22 16.433 73.276 16.633 ;
 RECT 72.38 16.433 72.436 16.633 ;
 RECT 72.212 16.433 72.268 16.633 ;
 RECT 72.716 16.433 72.772 16.633 ;
 RECT 72.548 16.433 72.604 16.633 ;
 RECT 71.708 16.433 71.764 16.633 ;
 RECT 71.54 16.433 71.596 16.633 ;
 RECT 72.044 16.433 72.1 16.633 ;
 RECT 71.876 16.433 71.932 16.633 ;
 RECT 71.036 16.433 71.092 16.633 ;
 RECT 70.868 16.433 70.924 16.633 ;
 RECT 71.372 16.433 71.428 16.633 ;
 RECT 71.204 16.433 71.26 16.633 ;
 RECT 70.364 16.433 70.42 16.633 ;
 RECT 70.7 16.433 70.756 16.633 ;
 RECT 70.532 16.433 70.588 16.633 ;
 RECT 74.396 17.2925 74.452 17.4925 ;
 RECT 74.228 17.2915 74.284 17.4915 ;
 RECT 74.732 17.106 74.788 17.306 ;
 RECT 74.564 17.2925 74.62 17.4925 ;
 RECT 73.724 17.2925 73.78 17.4925 ;
 RECT 73.556 17.2915 73.612 17.4915 ;
 RECT 74.06 17.106 74.116 17.306 ;
 RECT 73.892 17.2925 73.948 17.4925 ;
 RECT 73.052 17.2925 73.108 17.4925 ;
 RECT 72.884 17.2915 72.94 17.4915 ;
 RECT 73.388 17.106 73.444 17.306 ;
 RECT 73.22 17.2925 73.276 17.4925 ;
 RECT 72.38 17.2925 72.436 17.4925 ;
 RECT 72.212 17.2915 72.268 17.4915 ;
 RECT 72.716 17.106 72.772 17.306 ;
 RECT 72.548 17.2925 72.604 17.4925 ;
 RECT 71.708 17.2925 71.764 17.4925 ;
 RECT 71.54 17.2915 71.596 17.4915 ;
 RECT 72.044 17.106 72.1 17.306 ;
 RECT 71.876 17.2925 71.932 17.4925 ;
 RECT 71.036 17.2925 71.092 17.4925 ;
 RECT 70.868 17.2915 70.924 17.4915 ;
 RECT 71.372 17.106 71.428 17.306 ;
 RECT 71.204 17.2925 71.26 17.4925 ;
 RECT 70.364 17.2925 70.42 17.4925 ;
 RECT 70.7 17.106 70.756 17.306 ;
 RECT 70.532 17.2925 70.588 17.4925 ;
 END
 END vccdgt_1p0.gds1271
 PIN vccdgt_1p0.gds1272
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 24.383 0.654 24.583 ;
 END
 END vccdgt_1p0.gds1272
 PIN vccdgt_1p0.gds1273
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 23.123 0.654 23.323 ;
 END
 END vccdgt_1p0.gds1273
 PIN vccdgt_1p0.gds1274
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 21.863 0.654 22.063 ;
 END
 END vccdgt_1p0.gds1274
 PIN vccdgt_1p0.gds1275
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 20.603 0.654 20.803 ;
 END
 END vccdgt_1p0.gds1275
 PIN vccdgt_1p0.gds1276
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.454 23.138 0.494 23.338 ;
 END
 END vccdgt_1p0.gds1276
 PIN vccdgt_1p0.gds1277
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.566 23.357 1.622 23.557 ;
 END
 END vccdgt_1p0.gds1277
 PIN vccdgt_1p0.gds1278
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.742 23.0845 0.788 23.2845 ;
 END
 END vccdgt_1p0.gds1278
 PIN vccdgt_1p0.gds1279
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.114 23.037 1.154 23.237 ;
 END
 END vccdgt_1p0.gds1279
 PIN vccdgt_1p0.gds1280
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.966 23.1265 1.026 23.3265 ;
 END
 END vccdgt_1p0.gds1280
 PIN vccdgt_1p0.gds1281
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.986 23.0765 2.042 23.2765 ;
 END
 END vccdgt_1p0.gds1281
 PIN vccdgt_1p0.gds1282
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.69 20.6635 3.73 20.8635 ;
 END
 END vccdgt_1p0.gds1282
 PIN vccdgt_1p0.gds1283
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.326 23.1185 2.382 23.3185 ;
 END
 END vccdgt_1p0.gds1283
 PIN vccdgt_1p0.gds1284
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.806 23.086 1.882 23.286 ;
 END
 END vccdgt_1p0.gds1284
 PIN vccdgt_1p0.gds1285
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.882 21.034 3.922 21.234 ;
 END
 END vccdgt_1p0.gds1285
 PIN vccdgt_1p0.gds1286
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.646 23.0785 2.722 23.2785 ;
 END
 END vccdgt_1p0.gds1286
 PIN vccdgt_1p0.gds1287
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.098 25.3395 5.138 25.5395 ;
 END
 END vccdgt_1p0.gds1287
 PIN vccdgt_1p0.gds1288
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.634 23.047 4.674 23.247 ;
 END
 END vccdgt_1p0.gds1288
 PIN vccdgt_1p0.gds1289
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.478 23.014 3.538 23.214 ;
 END
 END vccdgt_1p0.gds1289
 PIN vccdgt_1p0.gds1290
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.09 25.3945 4.13 25.5945 ;
 END
 END vccdgt_1p0.gds1290
 PIN vccdgt_1p0.gds1291
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.906 25.186 4.946 25.386 ;
 END
 END vccdgt_1p0.gds1291
 PIN vccdgt_1p0.gds1292
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.362 23.022 4.418 23.222 ;
 END
 END vccdgt_1p0.gds1292
 PIN vccdgt_1p0.gds1293
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.762 23.138 4.818 23.338 ;
 END
 END vccdgt_1p0.gds1293
 PIN vccdgt_1p0.gds1294
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.486 23.002 2.542 23.202 ;
 END
 END vccdgt_1p0.gds1294
 PIN vccdgt_1p0.gds1295
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 1.232 20.88 1.288 21.08 ;
 RECT 1.568 20.895 1.624 21.095 ;
 RECT 1.82 20.895 1.876 21.095 ;
 RECT 2.072 21.009 2.128 21.189 ;
 RECT 2.492 20.5085 2.548 20.7085 ;
 RECT 2.996 21.007 3.052 21.189 ;
 RECT 3.164 21.007 3.22 21.183 ;
 RECT 1.232 22.14 1.288 22.34 ;
 RECT 1.568 22.155 1.624 22.355 ;
 RECT 1.82 22.155 1.876 22.355 ;
 RECT 2.072 22.269 2.128 22.449 ;
 RECT 2.996 22.267 3.052 22.449 ;
 RECT 3.164 22.267 3.22 22.443 ;
 RECT 2.492 21.7685 2.548 21.9685 ;
 RECT 1.232 23.4 1.288 23.6 ;
 RECT 1.568 23.415 1.624 23.615 ;
 RECT 1.82 23.415 1.876 23.615 ;
 RECT 2.072 23.529 2.128 23.709 ;
 RECT 2.996 23.527 3.052 23.709 ;
 RECT 3.164 23.527 3.22 23.703 ;
 RECT 2.492 23.0285 2.548 23.2285 ;
 RECT 1.232 24.66 1.288 24.86 ;
 RECT 1.568 24.675 1.624 24.875 ;
 RECT 1.82 24.675 1.876 24.875 ;
 RECT 2.072 24.789 2.128 24.969 ;
 RECT 2.996 24.787 3.052 24.969 ;
 RECT 3.164 24.787 3.22 24.963 ;
 RECT 2.492 24.2885 2.548 24.4885 ;
 RECT 0.812 20.913 0.868 21.113 ;
 RECT 0.644 20.913 0.7 21.113 ;
 RECT 0.98 20.913 1.036 21.113 ;
 RECT 0.812 22.173 0.868 22.373 ;
 RECT 0.644 22.173 0.7 22.373 ;
 RECT 0.98 22.173 1.036 22.373 ;
 RECT 0.812 23.433 0.868 23.633 ;
 RECT 0.644 23.433 0.7 23.633 ;
 RECT 0.98 23.433 1.036 23.633 ;
 RECT 0.812 24.693 0.868 24.893 ;
 RECT 0.644 24.693 0.7 24.893 ;
 RECT 0.98 24.693 1.036 24.893 ;
 RECT 4.088 24.2375 4.144 24.4375 ;
 RECT 4.676 24.2375 4.732 24.4375 ;
 RECT 4.424 24.2375 4.48 24.4375 ;
 RECT 5.012 24.2375 5.068 24.4375 ;
 RECT 4.844 24.2375 4.9 24.4375 ;
 RECT 4.088 22.9775 4.144 23.1775 ;
 RECT 4.676 22.9775 4.732 23.1775 ;
 RECT 4.424 22.9775 4.48 23.1775 ;
 RECT 5.012 22.9775 5.068 23.1775 ;
 RECT 4.844 22.9775 4.9 23.1775 ;
 RECT 4.088 21.7175 4.144 21.9175 ;
 RECT 4.676 21.7175 4.732 21.9175 ;
 RECT 4.424 21.7175 4.48 21.9175 ;
 RECT 5.012 21.7175 5.068 21.9175 ;
 RECT 4.844 21.7175 4.9 21.9175 ;
 RECT 4.088 20.4575 4.144 20.6575 ;
 RECT 4.676 20.4575 4.732 20.6575 ;
 RECT 4.424 20.4575 4.48 20.6575 ;
 RECT 5.012 20.4575 5.068 20.6575 ;
 RECT 4.844 20.4575 4.9 20.6575 ;
 END
 END vccdgt_1p0.gds1295
 PIN vccdgt_1p0.gds1296
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.626 23.644 5.666 23.844 ;
 END
 END vccdgt_1p0.gds1296
 PIN vccdgt_1p0.gds1297
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.33 23.873 6.37 24.073 ;
 END
 END vccdgt_1p0.gds1297
 PIN vccdgt_1p0.gds1298
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.862 23.0165 6.918 23.2165 ;
 END
 END vccdgt_1p0.gds1298
 PIN vccdgt_1p0.gds1299
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.074 23.026 6.114 23.226 ;
 END
 END vccdgt_1p0.gds1299
 PIN vccdgt_1p0.gds1300
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.306 23.0165 5.346 23.2165 ;
 END
 END vccdgt_1p0.gds1300
 PIN vccdgt_1p0.gds1301
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.818 22.9795 5.858 23.1795 ;
 END
 END vccdgt_1p0.gds1301
 PIN vccdgt_1p0.gds1302
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.498 24.875 5.538 25.075 ;
 END
 END vccdgt_1p0.gds1302
 PIN vccdgt_1p0.gds1303
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.202 23.0935 6.242 23.2935 ;
 END
 END vccdgt_1p0.gds1303
 PIN vccdgt_1p0.gds1304
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.67 23.033 6.71 23.233 ;
 END
 END vccdgt_1p0.gds1304
 PIN vccdgt_1p0.gds1305
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.348 24.2885 5.404 24.4885 ;
 RECT 6.02 24.2375 6.076 24.4375 ;
 RECT 5.684 24.3165 5.74 24.5165 ;
 RECT 6.356 24.3165 6.412 24.5165 ;
 RECT 5.348 23.0285 5.404 23.2285 ;
 RECT 6.02 22.9775 6.076 23.1775 ;
 RECT 5.684 23.0565 5.74 23.2565 ;
 RECT 6.356 23.0565 6.412 23.2565 ;
 RECT 5.348 21.7685 5.404 21.9685 ;
 RECT 6.02 21.7175 6.076 21.9175 ;
 RECT 5.684 21.7965 5.74 21.9965 ;
 RECT 6.356 21.7965 6.412 21.9965 ;
 RECT 6.02 20.4575 6.076 20.6575 ;
 RECT 5.348 20.5085 5.404 20.7085 ;
 RECT 5.684 20.5365 5.74 20.7365 ;
 RECT 6.356 20.5365 6.412 20.7365 ;
 END
 END vccdgt_1p0.gds1305
 PIN vccdgt_1p0.gds1306
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.522 22.5115 14.578 22.7115 ;
 END
 END vccdgt_1p0.gds1306
 PIN vccdgt_1p0.gds1307
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.342 23.5335 13.398 23.7335 ;
 END
 END vccdgt_1p0.gds1307
 PIN vccdgt_1p0.gds1308
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.186 24.033 15.226 24.233 ;
 END
 END vccdgt_1p0.gds1308
 PIN vccdgt_1p0.gds1309
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.182 23.914 14.238 24.114 ;
 END
 END vccdgt_1p0.gds1309
 PIN vccdgt_1p0.gds1310
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.502 23.904 13.558 24.104 ;
 END
 END vccdgt_1p0.gds1310
 PIN vccdgt_1p0.gds1311
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.162 23.103 13.238 23.303 ;
 END
 END vccdgt_1p0.gds1311
 PIN vccdgt_1p0.gds1312
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.766 22.773 14.806 22.973 ;
 END
 END vccdgt_1p0.gds1312
 PIN vccdgt_1p0.gds1313
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.002 23.914 14.078 24.114 ;
 END
 END vccdgt_1p0.gds1313
 PIN vccdgt_1p0.gds1314
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.958 24.0415 14.998 24.2415 ;
 END
 END vccdgt_1p0.gds1314
 PIN vccdgt_1p0.gds1315
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.678 23.4525 12.718 23.6525 ;
 END
 END vccdgt_1p0.gds1315
 PIN vccdgt_1p0.gds1316
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.402 23.0785 12.462 23.2785 ;
 END
 END vccdgt_1p0.gds1316
 PIN vccdgt_1p0.gds1317
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 14.756 21.677 14.812 21.877 ;
 RECT 14.756 22.937 14.812 23.137 ;
 RECT 14.756 24.197 14.812 24.397 ;
 RECT 14 25.34 14.056 25.54 ;
 RECT 14 21.56 14.056 21.76 ;
 RECT 14 22.82 14.056 23.02 ;
 RECT 14 24.08 14.056 24.28 ;
 RECT 14.924 25.024 14.98 25.224 ;
 RECT 14.42 25.444 14.476 25.644 ;
 RECT 14.924 23.764 14.98 23.964 ;
 RECT 14.588 24.197 14.644 24.397 ;
 RECT 14.42 24.184 14.476 24.384 ;
 RECT 14.924 22.504 14.98 22.704 ;
 RECT 14.588 22.937 14.644 23.137 ;
 RECT 14.42 22.924 14.476 23.124 ;
 RECT 14.924 21.244 14.98 21.444 ;
 RECT 14.588 21.677 14.644 21.877 ;
 RECT 14.42 21.664 14.476 21.864 ;
 END
 END vccdgt_1p0.gds1317
 PIN vccdgt_1p0.gds1318
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 20.926 16.57 21.126 ;
 END
 END vccdgt_1p0.gds1318
 PIN vccdgt_1p0.gds1319
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 22.186 16.57 22.386 ;
 END
 END vccdgt_1p0.gds1319
 PIN vccdgt_1p0.gds1320
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 23.446 16.57 23.646 ;
 END
 END vccdgt_1p0.gds1320
 PIN vccdgt_1p0.gds1321
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 24.706 16.57 24.906 ;
 END
 END vccdgt_1p0.gds1321
 PIN vccdgt_1p0.gds1322
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.866 23.7715 15.926 23.9715 ;
 END
 END vccdgt_1p0.gds1322
 PIN vccdgt_1p0.gds1323
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.838 24.7935 16.894 24.9935 ;
 END
 END vccdgt_1p0.gds1323
 PIN vccdgt_1p0.gds1324
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.674 24.1635 16.734 24.3635 ;
 END
 END vccdgt_1p0.gds1324
 PIN vccdgt_1p0.gds1325
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.018 24.786 17.074 24.986 ;
 END
 END vccdgt_1p0.gds1325
 PIN vccdgt_1p0.gds1326
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.03 23.929 16.076 24.129 ;
 END
 END vccdgt_1p0.gds1326
 PIN vccdgt_1p0.gds1327
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.314 23.1415 15.354 23.3415 ;
 END
 END vccdgt_1p0.gds1327
 PIN vccdgt_1p0.gds1328
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.338 23.2185 17.414 23.4185 ;
 END
 END vccdgt_1p0.gds1328
 PIN vccdgt_1p0.gds1329
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.114 23.0785 18.174 23.2785 ;
 END
 END vccdgt_1p0.gds1329
 PIN vccdgt_1p0.gds1330
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.858 24.73 17.898 24.93 ;
 END
 END vccdgt_1p0.gds1330
 PIN vccdgt_1p0.gds1331
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.522 22.8605 15.582 23.0605 ;
 END
 END vccdgt_1p0.gds1331
 PIN vccdgt_1p0.gds1332
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.598 22.6645 17.654 22.8645 ;
 END
 END vccdgt_1p0.gds1332
 PIN vccdgt_1p0.gds1333
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.178 23.05 17.234 23.25 ;
 END
 END vccdgt_1p0.gds1333
 PIN vccdgt_1p0.gds1334
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 15.932 20.48 15.988 20.68 ;
 RECT 15.932 21.74 15.988 21.94 ;
 RECT 15.932 23 15.988 23.2 ;
 RECT 15.932 24.26 15.988 24.46 ;
 RECT 15.764 25.1 15.82 25.3 ;
 RECT 15.512 25.352 15.568 25.552 ;
 RECT 15.26 25.439 15.316 25.639 ;
 RECT 15.764 23.84 15.82 24.04 ;
 RECT 15.512 24.092 15.568 24.292 ;
 RECT 15.26 24.179 15.316 24.379 ;
 RECT 16.1 24.197 16.156 24.397 ;
 RECT 15.764 22.58 15.82 22.78 ;
 RECT 15.512 22.832 15.568 23.032 ;
 RECT 15.26 22.919 15.316 23.119 ;
 RECT 16.1 22.937 16.156 23.137 ;
 RECT 15.764 21.32 15.82 21.52 ;
 RECT 15.512 21.572 15.568 21.772 ;
 RECT 15.26 21.659 15.316 21.859 ;
 RECT 16.1 21.677 16.156 21.877 ;
 END
 END vccdgt_1p0.gds1334
 PIN vccdgt_1p0.gds1335
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.93 23.138 23.97 23.338 ;
 END
 END vccdgt_1p0.gds1335
 PIN vccdgt_1p0.gds1336
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.658 22.923 23.698 23.123 ;
 END
 END vccdgt_1p0.gds1336
 PIN vccdgt_1p0.gds1337
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.214 23.103 30.29 23.303 ;
 END
 END vccdgt_1p0.gds1337
 PIN vccdgt_1p0.gds1338
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.73 23.4525 29.77 23.6525 ;
 END
 END vccdgt_1p0.gds1338
 PIN vccdgt_1p0.gds1339
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.454 23.0785 29.514 23.2785 ;
 END
 END vccdgt_1p0.gds1339
 PIN vccdgt_1p0.gds1340
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 20.926 33.622 21.126 ;
 END
 END vccdgt_1p0.gds1340
 PIN vccdgt_1p0.gds1341
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 22.186 33.622 22.386 ;
 END
 END vccdgt_1p0.gds1341
 PIN vccdgt_1p0.gds1342
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 24.706 33.622 24.906 ;
 END
 END vccdgt_1p0.gds1342
 PIN vccdgt_1p0.gds1343
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 23.446 33.622 23.646 ;
 END
 END vccdgt_1p0.gds1343
 PIN vccdgt_1p0.gds1344
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.574 22.5115 31.63 22.7115 ;
 END
 END vccdgt_1p0.gds1344
 PIN vccdgt_1p0.gds1345
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.918 23.7715 32.978 23.9715 ;
 END
 END vccdgt_1p0.gds1345
 PIN vccdgt_1p0.gds1346
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.238 23.7715 32.278 23.9715 ;
 END
 END vccdgt_1p0.gds1346
 PIN vccdgt_1p0.gds1347
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.394 23.5335 30.45 23.7335 ;
 END
 END vccdgt_1p0.gds1347
 PIN vccdgt_1p0.gds1348
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.89 24.7935 33.946 24.9935 ;
 END
 END vccdgt_1p0.gds1348
 PIN vccdgt_1p0.gds1349
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.726 24.1635 33.786 24.3635 ;
 END
 END vccdgt_1p0.gds1349
 PIN vccdgt_1p0.gds1350
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.07 24.786 34.126 24.986 ;
 END
 END vccdgt_1p0.gds1350
 PIN vccdgt_1p0.gds1351
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.39 23.2185 34.466 23.4185 ;
 END
 END vccdgt_1p0.gds1351
 PIN vccdgt_1p0.gds1352
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.082 23.929 33.128 24.129 ;
 END
 END vccdgt_1p0.gds1352
 PIN vccdgt_1p0.gds1353
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.366 23.718 32.406 23.918 ;
 END
 END vccdgt_1p0.gds1353
 PIN vccdgt_1p0.gds1354
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.554 23.904 30.61 24.104 ;
 END
 END vccdgt_1p0.gds1354
 PIN vccdgt_1p0.gds1355
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.818 22.773 31.858 22.973 ;
 END
 END vccdgt_1p0.gds1355
 PIN vccdgt_1p0.gds1356
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.234 23.914 31.29 24.114 ;
 END
 END vccdgt_1p0.gds1356
 PIN vccdgt_1p0.gds1357
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.91 24.73 34.95 24.93 ;
 END
 END vccdgt_1p0.gds1357
 PIN vccdgt_1p0.gds1358
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.574 22.8605 32.634 23.0605 ;
 END
 END vccdgt_1p0.gds1358
 PIN vccdgt_1p0.gds1359
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.65 22.6645 34.706 22.8645 ;
 END
 END vccdgt_1p0.gds1359
 PIN vccdgt_1p0.gds1360
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.01 24.0415 32.05 24.2415 ;
 END
 END vccdgt_1p0.gds1360
 PIN vccdgt_1p0.gds1361
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.166 23.0785 35.226 23.2785 ;
 END
 END vccdgt_1p0.gds1361
 PIN vccdgt_1p0.gds1362
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.054 23.914 31.13 24.114 ;
 END
 END vccdgt_1p0.gds1362
 PIN vccdgt_1p0.gds1363
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.23 23.05 34.286 23.25 ;
 END
 END vccdgt_1p0.gds1363
 PIN vccdgt_1p0.gds1364
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 33.152 21.677 33.208 21.877 ;
 RECT 31.052 22.82 31.108 23.02 ;
 RECT 31.808 22.937 31.864 23.137 ;
 RECT 33.152 24.197 33.208 24.397 ;
 RECT 31.052 25.34 31.108 25.54 ;
 RECT 31.976 25.024 32.032 25.224 ;
 RECT 32.816 25.1 32.872 25.3 ;
 RECT 32.564 25.352 32.62 25.552 ;
 RECT 31.472 25.444 31.528 25.644 ;
 RECT 32.312 25.439 32.368 25.639 ;
 RECT 31.052 24.08 31.108 24.28 ;
 RECT 31.808 24.197 31.864 24.397 ;
 RECT 32.984 24.26 33.04 24.46 ;
 RECT 31.976 23.764 32.032 23.964 ;
 RECT 32.816 23.84 32.872 24.04 ;
 RECT 32.564 24.092 32.62 24.292 ;
 RECT 32.312 24.179 32.368 24.379 ;
 RECT 31.64 24.197 31.696 24.397 ;
 RECT 31.472 24.184 31.528 24.384 ;
 RECT 31.976 22.504 32.032 22.704 ;
 RECT 32.816 22.58 32.872 22.78 ;
 RECT 32.564 22.832 32.62 23.032 ;
 RECT 32.984 23 33.04 23.2 ;
 RECT 31.64 22.937 31.696 23.137 ;
 RECT 33.152 22.937 33.208 23.137 ;
 RECT 31.472 22.924 31.528 23.124 ;
 RECT 32.312 22.919 32.368 23.119 ;
 RECT 31.052 21.56 31.108 21.76 ;
 RECT 31.808 21.677 31.864 21.877 ;
 RECT 32.984 21.74 33.04 21.94 ;
 RECT 31.976 21.244 32.032 21.444 ;
 RECT 32.816 21.32 32.872 21.52 ;
 RECT 32.564 21.572 32.62 21.772 ;
 RECT 32.312 21.659 32.368 21.859 ;
 RECT 31.64 21.677 31.696 21.877 ;
 RECT 31.472 21.664 31.528 21.864 ;
 RECT 32.984 20.48 33.04 20.68 ;
 END
 END vccdgt_1p0.gds1364
 PIN vccdgt_1p0.gds1365
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.982 23.138 41.022 23.338 ;
 END
 END vccdgt_1p0.gds1365
 PIN vccdgt_1p0.gds1366
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.71 22.923 40.75 23.123 ;
 END
 END vccdgt_1p0.gds1366
 PIN vccdgt_1p0.gds1367
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.446 23.5335 47.502 23.7335 ;
 END
 END vccdgt_1p0.gds1367
 PIN vccdgt_1p0.gds1368
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.97 23.7715 50.03 23.9715 ;
 END
 END vccdgt_1p0.gds1368
 PIN vccdgt_1p0.gds1369
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.626 22.5115 48.682 22.7115 ;
 END
 END vccdgt_1p0.gds1369
 PIN vccdgt_1p0.gds1370
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.29 23.7715 49.33 23.9715 ;
 END
 END vccdgt_1p0.gds1370
 PIN vccdgt_1p0.gds1371
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.418 23.718 49.458 23.918 ;
 END
 END vccdgt_1p0.gds1371
 PIN vccdgt_1p0.gds1372
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.606 23.904 47.662 24.104 ;
 END
 END vccdgt_1p0.gds1372
 PIN vccdgt_1p0.gds1373
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.266 23.103 47.342 23.303 ;
 END
 END vccdgt_1p0.gds1373
 PIN vccdgt_1p0.gds1374
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.106 23.914 48.182 24.114 ;
 END
 END vccdgt_1p0.gds1374
 PIN vccdgt_1p0.gds1375
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.87 22.773 48.91 22.973 ;
 END
 END vccdgt_1p0.gds1375
 PIN vccdgt_1p0.gds1376
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.286 23.914 48.342 24.114 ;
 END
 END vccdgt_1p0.gds1376
 PIN vccdgt_1p0.gds1377
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.062 24.0415 49.102 24.2415 ;
 END
 END vccdgt_1p0.gds1377
 PIN vccdgt_1p0.gds1378
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.626 22.8605 49.686 23.0605 ;
 END
 END vccdgt_1p0.gds1378
 PIN vccdgt_1p0.gds1379
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.782 23.4525 46.822 23.6525 ;
 END
 END vccdgt_1p0.gds1379
 PIN vccdgt_1p0.gds1380
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.134 23.929 50.18 24.129 ;
 END
 END vccdgt_1p0.gds1380
 PIN vccdgt_1p0.gds1381
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.506 23.0785 46.566 23.2785 ;
 END
 END vccdgt_1p0.gds1381
 PIN vccdgt_1p0.gds1382
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 50.036 20.48 50.092 20.68 ;
 RECT 48.86 21.677 48.916 21.877 ;
 RECT 50.036 21.74 50.092 21.94 ;
 RECT 48.86 22.937 48.916 23.137 ;
 RECT 50.036 23 50.092 23.2 ;
 RECT 48.86 24.197 48.916 24.397 ;
 RECT 50.036 24.26 50.092 24.46 ;
 RECT 48.104 21.56 48.16 21.76 ;
 RECT 48.104 22.82 48.16 23.02 ;
 RECT 48.104 24.08 48.16 24.28 ;
 RECT 48.104 25.34 48.16 25.54 ;
 RECT 49.028 25.024 49.084 25.224 ;
 RECT 49.868 25.1 49.924 25.3 ;
 RECT 49.616 25.352 49.672 25.552 ;
 RECT 49.364 25.439 49.42 25.639 ;
 RECT 48.524 25.444 48.58 25.644 ;
 RECT 49.028 23.764 49.084 23.964 ;
 RECT 49.868 23.84 49.924 24.04 ;
 RECT 49.616 24.092 49.672 24.292 ;
 RECT 49.364 24.179 49.42 24.379 ;
 RECT 48.692 24.197 48.748 24.397 ;
 RECT 50.204 24.197 50.26 24.397 ;
 RECT 48.524 24.184 48.58 24.384 ;
 RECT 49.028 22.504 49.084 22.704 ;
 RECT 49.868 22.58 49.924 22.78 ;
 RECT 49.616 22.832 49.672 23.032 ;
 RECT 49.364 22.919 49.42 23.119 ;
 RECT 48.692 22.937 48.748 23.137 ;
 RECT 50.204 22.937 50.26 23.137 ;
 RECT 48.524 22.924 48.58 23.124 ;
 RECT 49.028 21.244 49.084 21.444 ;
 RECT 49.868 21.32 49.924 21.52 ;
 RECT 49.616 21.572 49.672 21.772 ;
 RECT 49.364 21.659 49.42 21.859 ;
 RECT 48.692 21.677 48.748 21.877 ;
 RECT 50.204 21.677 50.26 21.877 ;
 RECT 48.524 21.664 48.58 21.864 ;
 END
 END vccdgt_1p0.gds1382
 PIN vccdgt_1p0.gds1383
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 20.926 50.674 21.126 ;
 END
 END vccdgt_1p0.gds1383
 PIN vccdgt_1p0.gds1384
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 22.186 50.674 22.386 ;
 END
 END vccdgt_1p0.gds1384
 PIN vccdgt_1p0.gds1385
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 23.446 50.674 23.646 ;
 END
 END vccdgt_1p0.gds1385
 PIN vccdgt_1p0.gds1386
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 24.706 50.674 24.906 ;
 END
 END vccdgt_1p0.gds1386
 PIN vccdgt_1p0.gds1387
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.942 24.7935 50.998 24.9935 ;
 END
 END vccdgt_1p0.gds1387
 PIN vccdgt_1p0.gds1388
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.778 24.1635 50.838 24.3635 ;
 END
 END vccdgt_1p0.gds1388
 PIN vccdgt_1p0.gds1389
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.122 24.786 51.178 24.986 ;
 END
 END vccdgt_1p0.gds1389
 PIN vccdgt_1p0.gds1390
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.442 23.2185 51.518 23.4185 ;
 END
 END vccdgt_1p0.gds1390
 PIN vccdgt_1p0.gds1391
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.218 23.0785 52.278 23.2785 ;
 END
 END vccdgt_1p0.gds1391
 PIN vccdgt_1p0.gds1392
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.962 24.73 52.002 24.93 ;
 END
 END vccdgt_1p0.gds1392
 PIN vccdgt_1p0.gds1393
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.282 23.05 51.338 23.25 ;
 END
 END vccdgt_1p0.gds1393
 PIN vccdgt_1p0.gds1394
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.702 22.6645 51.758 22.8645 ;
 END
 END vccdgt_1p0.gds1394
 PIN vccdgt_1p0.gds1395
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.034 23.138 58.074 23.338 ;
 END
 END vccdgt_1p0.gds1395
 PIN vccdgt_1p0.gds1396
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.762 22.923 57.802 23.123 ;
 END
 END vccdgt_1p0.gds1396
 PIN vccdgt_1p0.gds1397
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.498 23.5335 64.554 23.7335 ;
 END
 END vccdgt_1p0.gds1397
 PIN vccdgt_1p0.gds1398
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.658 23.904 64.714 24.104 ;
 END
 END vccdgt_1p0.gds1398
 PIN vccdgt_1p0.gds1399
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.318 23.103 64.394 23.303 ;
 END
 END vccdgt_1p0.gds1399
 PIN vccdgt_1p0.gds1400
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.834 23.4525 63.874 23.6525 ;
 END
 END vccdgt_1p0.gds1400
 PIN vccdgt_1p0.gds1401
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.158 23.914 65.234 24.114 ;
 END
 END vccdgt_1p0.gds1401
 PIN vccdgt_1p0.gds1402
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.558 23.0785 63.618 23.2785 ;
 END
 END vccdgt_1p0.gds1402
 PIN vccdgt_1p0.gds1403
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 65.156 25.34 65.212 25.54 ;
 RECT 65.156 24.08 65.212 24.28 ;
 RECT 65.156 22.82 65.212 23.02 ;
 RECT 65.156 21.56 65.212 21.76 ;
 END
 END vccdgt_1p0.gds1403
 PIN vccdgt_1p0.gds1404
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 23.446 67.726 23.646 ;
 END
 END vccdgt_1p0.gds1404
 PIN vccdgt_1p0.gds1405
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 24.706 67.726 24.906 ;
 END
 END vccdgt_1p0.gds1405
 PIN vccdgt_1p0.gds1406
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 22.186 67.726 22.386 ;
 END
 END vccdgt_1p0.gds1406
 PIN vccdgt_1p0.gds1407
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 20.926 67.726 21.126 ;
 END
 END vccdgt_1p0.gds1407
 PIN vccdgt_1p0.gds1408
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.678 22.5115 65.734 22.7115 ;
 END
 END vccdgt_1p0.gds1408
 PIN vccdgt_1p0.gds1409
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.022 23.7715 67.082 23.9715 ;
 END
 END vccdgt_1p0.gds1409
 PIN vccdgt_1p0.gds1410
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.342 23.7715 66.382 23.9715 ;
 END
 END vccdgt_1p0.gds1410
 PIN vccdgt_1p0.gds1411
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.994 24.7935 68.05 24.9935 ;
 END
 END vccdgt_1p0.gds1411
 PIN vccdgt_1p0.gds1412
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.83 24.1635 67.89 24.3635 ;
 END
 END vccdgt_1p0.gds1412
 PIN vccdgt_1p0.gds1413
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.174 24.786 68.23 24.986 ;
 END
 END vccdgt_1p0.gds1413
 PIN vccdgt_1p0.gds1414
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.494 23.2185 68.57 23.4185 ;
 END
 END vccdgt_1p0.gds1414
 PIN vccdgt_1p0.gds1415
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.47 23.718 66.51 23.918 ;
 END
 END vccdgt_1p0.gds1415
 PIN vccdgt_1p0.gds1416
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.922 22.773 65.962 22.973 ;
 END
 END vccdgt_1p0.gds1416
 PIN vccdgt_1p0.gds1417
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.338 23.914 65.394 24.114 ;
 END
 END vccdgt_1p0.gds1417
 PIN vccdgt_1p0.gds1418
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.27 23.0785 69.33 23.2785 ;
 END
 END vccdgt_1p0.gds1418
 PIN vccdgt_1p0.gds1419
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.014 24.73 69.054 24.93 ;
 END
 END vccdgt_1p0.gds1419
 PIN vccdgt_1p0.gds1420
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.334 23.05 68.39 23.25 ;
 END
 END vccdgt_1p0.gds1420
 PIN vccdgt_1p0.gds1421
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.114 24.0415 66.154 24.2415 ;
 END
 END vccdgt_1p0.gds1421
 PIN vccdgt_1p0.gds1422
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.754 22.6645 68.81 22.8645 ;
 END
 END vccdgt_1p0.gds1422
 PIN vccdgt_1p0.gds1423
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.678 22.8605 66.738 23.0605 ;
 END
 END vccdgt_1p0.gds1423
 PIN vccdgt_1p0.gds1424
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.186 23.929 67.232 24.129 ;
 END
 END vccdgt_1p0.gds1424
 PIN vccdgt_1p0.gds1425
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 67.088 20.48 67.144 20.68 ;
 RECT 65.912 21.677 65.968 21.877 ;
 RECT 67.088 21.74 67.144 21.94 ;
 RECT 65.912 22.937 65.968 23.137 ;
 RECT 67.088 23 67.144 23.2 ;
 RECT 65.912 24.197 65.968 24.397 ;
 RECT 67.088 24.26 67.144 24.46 ;
 RECT 66.08 25.024 66.136 25.224 ;
 RECT 66.92 25.1 66.976 25.3 ;
 RECT 66.668 25.352 66.724 25.552 ;
 RECT 66.416 25.439 66.472 25.639 ;
 RECT 65.576 25.444 65.632 25.644 ;
 RECT 66.08 23.764 66.136 23.964 ;
 RECT 66.92 23.84 66.976 24.04 ;
 RECT 66.668 24.092 66.724 24.292 ;
 RECT 66.416 24.179 66.472 24.379 ;
 RECT 65.744 24.197 65.8 24.397 ;
 RECT 67.256 24.197 67.312 24.397 ;
 RECT 65.576 24.184 65.632 24.384 ;
 RECT 66.08 22.504 66.136 22.704 ;
 RECT 66.92 22.58 66.976 22.78 ;
 RECT 66.668 22.832 66.724 23.032 ;
 RECT 66.416 22.919 66.472 23.119 ;
 RECT 65.744 22.937 65.8 23.137 ;
 RECT 67.256 22.937 67.312 23.137 ;
 RECT 65.576 22.924 65.632 23.124 ;
 RECT 66.08 21.244 66.136 21.444 ;
 RECT 66.92 21.32 66.976 21.52 ;
 RECT 66.668 21.572 66.724 21.772 ;
 RECT 66.416 21.659 66.472 21.859 ;
 RECT 65.744 21.677 65.8 21.877 ;
 RECT 67.256 21.677 67.312 21.877 ;
 RECT 65.576 21.664 65.632 21.864 ;
 END
 END vccdgt_1p0.gds1425
 PIN vccdgt_1p0.gds1426
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 28.163 0.654 28.363 ;
 END
 END vccdgt_1p0.gds1426
 PIN vccdgt_1p0.gds1427
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 25.643 0.654 25.843 ;
 END
 END vccdgt_1p0.gds1427
 PIN vccdgt_1p0.gds1428
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.626 26.903 0.654 27.103 ;
 END
 END vccdgt_1p0.gds1428
 PIN vccdgt_1p0.gds1429
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.454 27.163 0.494 27.363 ;
 END
 END vccdgt_1p0.gds1429
 PIN vccdgt_1p0.gds1430
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.566 27.2405 1.622 27.4405 ;
 END
 END vccdgt_1p0.gds1430
 PIN vccdgt_1p0.gds1431
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.742 27.1755 0.788 27.3755 ;
 END
 END vccdgt_1p0.gds1431
 PIN vccdgt_1p0.gds1432
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.114 27.1565 1.154 27.3565 ;
 END
 END vccdgt_1p0.gds1432
 PIN vccdgt_1p0.gds1433
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.966 27.1585 1.026 27.3585 ;
 END
 END vccdgt_1p0.gds1433
 PIN vccdgt_1p0.gds1434
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.986 27.182 2.042 27.382 ;
 END
 END vccdgt_1p0.gds1434
 PIN vccdgt_1p0.gds1435
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.69 28.484 3.73 28.684 ;
 END
 END vccdgt_1p0.gds1435
 PIN vccdgt_1p0.gds1436
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.69 25.613 3.73 25.813 ;
 END
 END vccdgt_1p0.gds1436
 PIN vccdgt_1p0.gds1437
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.326 27.175 2.382 27.375 ;
 END
 END vccdgt_1p0.gds1437
 PIN vccdgt_1p0.gds1438
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.806 27.175 1.882 27.375 ;
 END
 END vccdgt_1p0.gds1438
 PIN vccdgt_1p0.gds1439
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.882 28.5475 3.922 28.7475 ;
 END
 END vccdgt_1p0.gds1439
 PIN vccdgt_1p0.gds1440
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.882 25.987 3.922 26.187 ;
 END
 END vccdgt_1p0.gds1440
 PIN vccdgt_1p0.gds1441
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.166 28.3555 3.206 28.5555 ;
 END
 END vccdgt_1p0.gds1441
 PIN vccdgt_1p0.gds1442
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.166 25.52 3.206 25.72 ;
 END
 END vccdgt_1p0.gds1442
 PIN vccdgt_1p0.gds1443
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.646 27.142 2.722 27.342 ;
 END
 END vccdgt_1p0.gds1443
 PIN vccdgt_1p0.gds1444
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.098 28.285 5.138 28.485 ;
 END
 END vccdgt_1p0.gds1444
 PIN vccdgt_1p0.gds1445
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.634 27.2045 4.674 27.4045 ;
 END
 END vccdgt_1p0.gds1445
 PIN vccdgt_1p0.gds1446
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.478 27.1225 3.538 27.3225 ;
 END
 END vccdgt_1p0.gds1446
 PIN vccdgt_1p0.gds1447
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.09 28.3675 4.13 28.5675 ;
 END
 END vccdgt_1p0.gds1447
 PIN vccdgt_1p0.gds1448
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.906 28.2585 4.946 28.4585 ;
 END
 END vccdgt_1p0.gds1448
 PIN vccdgt_1p0.gds1449
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.362 27.148 4.418 27.348 ;
 END
 END vccdgt_1p0.gds1449
 PIN vccdgt_1p0.gds1450
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.762 27.163 4.818 27.363 ;
 END
 END vccdgt_1p0.gds1450
 PIN vccdgt_1p0.gds1451
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.486 27.146 2.542 27.346 ;
 END
 END vccdgt_1p0.gds1451
 PIN vccdgt_1p0.gds1452
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 1.232 25.92 1.288 26.12 ;
 RECT 1.568 25.935 1.624 26.135 ;
 RECT 1.82 25.935 1.876 26.135 ;
 RECT 2.072 26.049 2.128 26.229 ;
 RECT 2.996 26.047 3.052 26.229 ;
 RECT 3.164 26.047 3.22 26.223 ;
 RECT 2.492 25.5485 2.548 25.7485 ;
 RECT 1.232 27.18 1.288 27.38 ;
 RECT 1.568 27.195 1.624 27.395 ;
 RECT 1.82 27.195 1.876 27.395 ;
 RECT 2.072 27.309 2.128 27.489 ;
 RECT 2.996 27.307 3.052 27.489 ;
 RECT 3.164 27.307 3.22 27.483 ;
 RECT 2.492 26.8085 2.548 27.0085 ;
 RECT 1.232 28.44 1.288 28.64 ;
 RECT 1.568 28.455 1.624 28.655 ;
 RECT 1.82 28.455 1.876 28.655 ;
 RECT 2.072 28.569 2.128 28.749 ;
 RECT 2.996 28.567 3.052 28.749 ;
 RECT 3.164 28.567 3.22 28.743 ;
 RECT 2.492 28.0685 2.548 28.2685 ;
 RECT 0.812 28.473 0.868 28.673 ;
 RECT 0.644 28.473 0.7 28.673 ;
 RECT 0.98 28.473 1.036 28.673 ;
 RECT 0.812 25.953 0.868 26.153 ;
 RECT 0.644 25.953 0.7 26.153 ;
 RECT 0.98 25.953 1.036 26.153 ;
 RECT 0.812 27.213 0.868 27.413 ;
 RECT 0.644 27.213 0.7 27.413 ;
 RECT 0.98 27.213 1.036 27.413 ;
 RECT 4.088 28.0175 4.144 28.2175 ;
 RECT 4.676 28.0175 4.732 28.2175 ;
 RECT 4.424 28.0175 4.48 28.2175 ;
 RECT 5.012 28.0175 5.068 28.2175 ;
 RECT 4.844 28.0175 4.9 28.2175 ;
 RECT 4.088 26.7575 4.144 26.9575 ;
 RECT 4.676 26.7575 4.732 26.9575 ;
 RECT 4.424 26.7575 4.48 26.9575 ;
 RECT 5.012 26.7575 5.068 26.9575 ;
 RECT 4.844 26.7575 4.9 26.9575 ;
 RECT 4.088 25.4975 4.144 25.6975 ;
 RECT 4.676 25.4975 4.732 25.6975 ;
 RECT 4.424 25.4975 4.48 25.6975 ;
 RECT 5.012 25.4975 5.068 25.6975 ;
 RECT 4.844 25.4975 4.9 25.6975 ;
 END
 END vccdgt_1p0.gds1452
 PIN vccdgt_1p0.gds1453
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.626 27.424 5.666 27.624 ;
 END
 END vccdgt_1p0.gds1453
 PIN vccdgt_1p0.gds1454
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.33 27.653 6.37 27.853 ;
 END
 END vccdgt_1p0.gds1454
 PIN vccdgt_1p0.gds1455
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.862 27.157 6.918 27.357 ;
 END
 END vccdgt_1p0.gds1455
 PIN vccdgt_1p0.gds1456
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.074 27.1645 6.114 27.3645 ;
 END
 END vccdgt_1p0.gds1456
 PIN vccdgt_1p0.gds1457
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.306 27.157 5.346 27.357 ;
 END
 END vccdgt_1p0.gds1457
 PIN vccdgt_1p0.gds1458
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.818 27.1325 5.858 27.3325 ;
 END
 END vccdgt_1p0.gds1458
 PIN vccdgt_1p0.gds1459
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.498 28.025 5.538 28.225 ;
 END
 END vccdgt_1p0.gds1459
 PIN vccdgt_1p0.gds1460
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.202 27.1915 6.242 27.3915 ;
 END
 END vccdgt_1p0.gds1460
 PIN vccdgt_1p0.gds1461
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.67 27.129 6.71 27.329 ;
 END
 END vccdgt_1p0.gds1461
 PIN vccdgt_1p0.gds1462
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.348 28.0685 5.404 28.2685 ;
 RECT 6.02 28.0175 6.076 28.2175 ;
 RECT 5.684 28.0965 5.74 28.2965 ;
 RECT 6.356 28.0965 6.412 28.2965 ;
 RECT 5.348 26.8085 5.404 27.0085 ;
 RECT 6.02 26.7575 6.076 26.9575 ;
 RECT 5.684 26.8365 5.74 27.0365 ;
 RECT 6.356 26.8365 6.412 27.0365 ;
 RECT 5.348 25.5485 5.404 25.7485 ;
 RECT 6.02 25.4975 6.076 25.6975 ;
 RECT 5.684 25.5765 5.74 25.7765 ;
 RECT 6.356 25.5765 6.412 25.7765 ;
 END
 END vccdgt_1p0.gds1462
 PIN vccdgt_1p0.gds1463
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.522 26.9215 14.578 27.1215 ;
 END
 END vccdgt_1p0.gds1463
 PIN vccdgt_1p0.gds1464
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.342 27.3135 13.398 27.5135 ;
 END
 END vccdgt_1p0.gds1464
 PIN vccdgt_1p0.gds1465
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.186 27.672 15.226 27.872 ;
 END
 END vccdgt_1p0.gds1465
 PIN vccdgt_1p0.gds1466
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.182 27.694 14.238 27.894 ;
 END
 END vccdgt_1p0.gds1466
 PIN vccdgt_1p0.gds1467
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.502 27.454 13.558 27.654 ;
 END
 END vccdgt_1p0.gds1467
 PIN vccdgt_1p0.gds1468
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.162 27.119 13.238 27.319 ;
 END
 END vccdgt_1p0.gds1468
 PIN vccdgt_1p0.gds1469
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.766 27.036 14.806 27.236 ;
 END
 END vccdgt_1p0.gds1469
 PIN vccdgt_1p0.gds1470
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.002 27.694 14.078 27.894 ;
 END
 END vccdgt_1p0.gds1470
 PIN vccdgt_1p0.gds1471
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.958 27.8215 14.998 28.0215 ;
 END
 END vccdgt_1p0.gds1471
 PIN vccdgt_1p0.gds1472
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.678 27.3475 12.718 27.5475 ;
 END
 END vccdgt_1p0.gds1472
 PIN vccdgt_1p0.gds1473
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.402 27.142 12.462 27.342 ;
 END
 END vccdgt_1p0.gds1473
 PIN vccdgt_1p0.gds1474
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 14.756 25.457 14.812 25.657 ;
 RECT 14.756 26.717 14.812 26.917 ;
 RECT 14.756 27.977 14.812 28.177 ;
 RECT 14 27.86 14.056 28.06 ;
 RECT 14 26.6 14.056 26.8 ;
 RECT 14.924 27.544 14.98 27.744 ;
 RECT 14.588 27.977 14.644 28.177 ;
 RECT 14.42 27.964 14.476 28.164 ;
 RECT 14.924 26.284 14.98 26.484 ;
 RECT 14.588 26.717 14.644 26.917 ;
 RECT 14.42 26.704 14.476 26.904 ;
 RECT 14.588 25.457 14.644 25.657 ;
 END
 END vccdgt_1p0.gds1474
 PIN vccdgt_1p0.gds1475
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 27.226 16.57 27.426 ;
 END
 END vccdgt_1p0.gds1475
 PIN vccdgt_1p0.gds1476
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 25.966 16.57 26.166 ;
 END
 END vccdgt_1p0.gds1476
 PIN vccdgt_1p0.gds1477
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.866 27.5515 15.926 27.7515 ;
 END
 END vccdgt_1p0.gds1477
 PIN vccdgt_1p0.gds1478
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 28.486 16.57 28.686 ;
 END
 END vccdgt_1p0.gds1478
 PIN vccdgt_1p0.gds1479
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.838 27.9435 16.894 28.1435 ;
 END
 END vccdgt_1p0.gds1479
 PIN vccdgt_1p0.gds1480
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.674 27.6025 16.734 27.8025 ;
 END
 END vccdgt_1p0.gds1480
 PIN vccdgt_1p0.gds1481
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.018 27.936 17.074 28.136 ;
 END
 END vccdgt_1p0.gds1481
 PIN vccdgt_1p0.gds1482
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.03 27.709 16.076 27.909 ;
 END
 END vccdgt_1p0.gds1482
 PIN vccdgt_1p0.gds1483
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.314 27.196 15.354 27.396 ;
 END
 END vccdgt_1p0.gds1483
 PIN vccdgt_1p0.gds1484
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.338 27.142 17.414 27.342 ;
 END
 END vccdgt_1p0.gds1484
 PIN vccdgt_1p0.gds1485
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.114 27.142 18.174 27.342 ;
 END
 END vccdgt_1p0.gds1485
 PIN vccdgt_1p0.gds1486
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.858 27.984 17.898 28.184 ;
 END
 END vccdgt_1p0.gds1486
 PIN vccdgt_1p0.gds1487
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.522 27.079 15.582 27.279 ;
 END
 END vccdgt_1p0.gds1487
 PIN vccdgt_1p0.gds1488
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.598 26.973 17.654 27.173 ;
 END
 END vccdgt_1p0.gds1488
 PIN vccdgt_1p0.gds1489
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.178 27.1435 17.234 27.3435 ;
 END
 END vccdgt_1p0.gds1489
 PIN vccdgt_1p0.gds1490
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 15.932 25.52 15.988 25.72 ;
 RECT 15.932 26.78 15.988 26.98 ;
 RECT 15.932 28.04 15.988 28.24 ;
 RECT 15.764 27.62 15.82 27.82 ;
 RECT 15.512 27.872 15.568 28.072 ;
 RECT 15.26 27.959 15.316 28.159 ;
 RECT 16.1 27.977 16.156 28.177 ;
 RECT 15.764 26.36 15.82 26.56 ;
 RECT 15.512 26.612 15.568 26.812 ;
 RECT 15.26 26.699 15.316 26.899 ;
 RECT 16.1 26.717 16.156 26.917 ;
 RECT 16.1 25.457 16.156 25.657 ;
 END
 END vccdgt_1p0.gds1490
 PIN vccdgt_1p0.gds1491
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.93 27.163 23.97 27.363 ;
 END
 END vccdgt_1p0.gds1491
 PIN vccdgt_1p0.gds1492
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.658 27.074 23.698 27.274 ;
 END
 END vccdgt_1p0.gds1492
 PIN vccdgt_1p0.gds1493
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.214 27.119 30.29 27.319 ;
 END
 END vccdgt_1p0.gds1493
 PIN vccdgt_1p0.gds1494
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.73 27.3475 29.77 27.5475 ;
 END
 END vccdgt_1p0.gds1494
 PIN vccdgt_1p0.gds1495
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.454 27.142 29.514 27.342 ;
 END
 END vccdgt_1p0.gds1495
 PIN vccdgt_1p0.gds1496
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 28.486 33.622 28.686 ;
 END
 END vccdgt_1p0.gds1496
 PIN vccdgt_1p0.gds1497
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 27.226 33.622 27.426 ;
 END
 END vccdgt_1p0.gds1497
 PIN vccdgt_1p0.gds1498
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 25.966 33.622 26.166 ;
 END
 END vccdgt_1p0.gds1498
 PIN vccdgt_1p0.gds1499
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.574 26.9215 31.63 27.1215 ;
 END
 END vccdgt_1p0.gds1499
 PIN vccdgt_1p0.gds1500
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.918 27.5515 32.978 27.7515 ;
 END
 END vccdgt_1p0.gds1500
 PIN vccdgt_1p0.gds1501
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.238 27.5515 32.278 27.7515 ;
 END
 END vccdgt_1p0.gds1501
 PIN vccdgt_1p0.gds1502
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.394 27.3135 30.45 27.5135 ;
 END
 END vccdgt_1p0.gds1502
 PIN vccdgt_1p0.gds1503
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.89 27.9435 33.946 28.1435 ;
 END
 END vccdgt_1p0.gds1503
 PIN vccdgt_1p0.gds1504
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.726 27.6025 33.786 27.8025 ;
 END
 END vccdgt_1p0.gds1504
 PIN vccdgt_1p0.gds1505
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.07 27.936 34.126 28.136 ;
 END
 END vccdgt_1p0.gds1505
 PIN vccdgt_1p0.gds1506
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.39 27.142 34.466 27.342 ;
 END
 END vccdgt_1p0.gds1506
 PIN vccdgt_1p0.gds1507
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.082 27.709 33.128 27.909 ;
 END
 END vccdgt_1p0.gds1507
 PIN vccdgt_1p0.gds1508
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.366 27.498 32.406 27.698 ;
 END
 END vccdgt_1p0.gds1508
 PIN vccdgt_1p0.gds1509
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.554 27.454 30.61 27.654 ;
 END
 END vccdgt_1p0.gds1509
 PIN vccdgt_1p0.gds1510
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.818 27.036 31.858 27.236 ;
 END
 END vccdgt_1p0.gds1510
 PIN vccdgt_1p0.gds1511
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.234 27.694 31.29 27.894 ;
 END
 END vccdgt_1p0.gds1511
 PIN vccdgt_1p0.gds1512
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.91 27.984 34.95 28.184 ;
 END
 END vccdgt_1p0.gds1512
 PIN vccdgt_1p0.gds1513
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.574 27.079 32.634 27.279 ;
 END
 END vccdgt_1p0.gds1513
 PIN vccdgt_1p0.gds1514
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.65 26.973 34.706 27.173 ;
 END
 END vccdgt_1p0.gds1514
 PIN vccdgt_1p0.gds1515
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.01 27.8215 32.05 28.0215 ;
 END
 END vccdgt_1p0.gds1515
 PIN vccdgt_1p0.gds1516
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.166 27.142 35.226 27.342 ;
 END
 END vccdgt_1p0.gds1516
 PIN vccdgt_1p0.gds1517
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.054 27.694 31.13 27.894 ;
 END
 END vccdgt_1p0.gds1517
 PIN vccdgt_1p0.gds1518
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.23 27.1435 34.286 27.3435 ;
 END
 END vccdgt_1p0.gds1518
 PIN vccdgt_1p0.gds1519
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 31.808 25.457 31.864 25.657 ;
 RECT 31.808 26.717 31.864 26.917 ;
 RECT 32.984 26.78 33.04 26.98 ;
 RECT 31.052 26.6 31.108 26.8 ;
 RECT 31.052 27.86 31.108 28.06 ;
 RECT 31.808 27.977 31.864 28.177 ;
 RECT 32.984 28.04 33.04 28.24 ;
 RECT 31.976 27.544 32.032 27.744 ;
 RECT 32.816 27.62 32.872 27.82 ;
 RECT 32.564 27.872 32.62 28.072 ;
 RECT 32.312 27.959 32.368 28.159 ;
 RECT 31.64 27.977 31.696 28.177 ;
 RECT 33.152 27.977 33.208 28.177 ;
 RECT 31.472 27.964 31.528 28.164 ;
 RECT 31.976 26.284 32.032 26.484 ;
 RECT 32.816 26.36 32.872 26.56 ;
 RECT 32.564 26.612 32.62 26.812 ;
 RECT 32.312 26.699 32.368 26.899 ;
 RECT 31.64 26.717 31.696 26.917 ;
 RECT 33.152 26.717 33.208 26.917 ;
 RECT 31.472 26.704 31.528 26.904 ;
 RECT 32.984 25.52 33.04 25.72 ;
 RECT 33.152 25.457 33.208 25.657 ;
 RECT 31.64 25.457 31.696 25.657 ;
 END
 END vccdgt_1p0.gds1519
 PIN vccdgt_1p0.gds1520
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.982 27.163 41.022 27.363 ;
 END
 END vccdgt_1p0.gds1520
 PIN vccdgt_1p0.gds1521
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.71 27.074 40.75 27.274 ;
 END
 END vccdgt_1p0.gds1521
 PIN vccdgt_1p0.gds1522
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.446 27.3135 47.502 27.5135 ;
 END
 END vccdgt_1p0.gds1522
 PIN vccdgt_1p0.gds1523
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.97 27.5515 50.03 27.7515 ;
 END
 END vccdgt_1p0.gds1523
 PIN vccdgt_1p0.gds1524
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.626 26.9215 48.682 27.1215 ;
 END
 END vccdgt_1p0.gds1524
 PIN vccdgt_1p0.gds1525
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.29 27.5515 49.33 27.7515 ;
 END
 END vccdgt_1p0.gds1525
 PIN vccdgt_1p0.gds1526
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.418 27.498 49.458 27.698 ;
 END
 END vccdgt_1p0.gds1526
 PIN vccdgt_1p0.gds1527
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.606 27.454 47.662 27.654 ;
 END
 END vccdgt_1p0.gds1527
 PIN vccdgt_1p0.gds1528
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.266 27.119 47.342 27.319 ;
 END
 END vccdgt_1p0.gds1528
 PIN vccdgt_1p0.gds1529
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.106 27.694 48.182 27.894 ;
 END
 END vccdgt_1p0.gds1529
 PIN vccdgt_1p0.gds1530
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.87 27.036 48.91 27.236 ;
 END
 END vccdgt_1p0.gds1530
 PIN vccdgt_1p0.gds1531
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.286 27.694 48.342 27.894 ;
 END
 END vccdgt_1p0.gds1531
 PIN vccdgt_1p0.gds1532
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.062 27.8215 49.102 28.0215 ;
 END
 END vccdgt_1p0.gds1532
 PIN vccdgt_1p0.gds1533
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.626 27.079 49.686 27.279 ;
 END
 END vccdgt_1p0.gds1533
 PIN vccdgt_1p0.gds1534
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.782 27.3475 46.822 27.5475 ;
 END
 END vccdgt_1p0.gds1534
 PIN vccdgt_1p0.gds1535
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.134 27.709 50.18 27.909 ;
 END
 END vccdgt_1p0.gds1535
 PIN vccdgt_1p0.gds1536
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.506 27.142 46.566 27.342 ;
 END
 END vccdgt_1p0.gds1536
 PIN vccdgt_1p0.gds1537
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 48.86 25.457 48.916 25.657 ;
 RECT 50.036 25.52 50.092 25.72 ;
 RECT 48.86 26.717 48.916 26.917 ;
 RECT 50.036 26.78 50.092 26.98 ;
 RECT 48.104 26.6 48.16 26.8 ;
 RECT 48.104 27.86 48.16 28.06 ;
 RECT 48.86 27.977 48.916 28.177 ;
 RECT 50.036 28.04 50.092 28.24 ;
 RECT 49.028 27.544 49.084 27.744 ;
 RECT 49.868 27.62 49.924 27.82 ;
 RECT 49.616 27.872 49.672 28.072 ;
 RECT 49.364 27.959 49.42 28.159 ;
 RECT 48.692 27.977 48.748 28.177 ;
 RECT 50.204 27.977 50.26 28.177 ;
 RECT 48.524 27.964 48.58 28.164 ;
 RECT 49.028 26.284 49.084 26.484 ;
 RECT 49.868 26.36 49.924 26.56 ;
 RECT 49.616 26.612 49.672 26.812 ;
 RECT 49.364 26.699 49.42 26.899 ;
 RECT 48.692 26.717 48.748 26.917 ;
 RECT 50.204 26.717 50.26 26.917 ;
 RECT 48.524 26.704 48.58 26.904 ;
 RECT 48.692 25.457 48.748 25.657 ;
 RECT 50.204 25.457 50.26 25.657 ;
 END
 END vccdgt_1p0.gds1537
 PIN vccdgt_1p0.gds1538
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 27.226 50.674 27.426 ;
 END
 END vccdgt_1p0.gds1538
 PIN vccdgt_1p0.gds1539
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 25.966 50.674 26.166 ;
 END
 END vccdgt_1p0.gds1539
 PIN vccdgt_1p0.gds1540
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 28.486 50.674 28.686 ;
 END
 END vccdgt_1p0.gds1540
 PIN vccdgt_1p0.gds1541
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.942 27.9435 50.998 28.1435 ;
 END
 END vccdgt_1p0.gds1541
 PIN vccdgt_1p0.gds1542
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.778 27.6025 50.838 27.8025 ;
 END
 END vccdgt_1p0.gds1542
 PIN vccdgt_1p0.gds1543
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.122 27.936 51.178 28.136 ;
 END
 END vccdgt_1p0.gds1543
 PIN vccdgt_1p0.gds1544
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.442 27.142 51.518 27.342 ;
 END
 END vccdgt_1p0.gds1544
 PIN vccdgt_1p0.gds1545
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.218 27.142 52.278 27.342 ;
 END
 END vccdgt_1p0.gds1545
 PIN vccdgt_1p0.gds1546
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.962 27.984 52.002 28.184 ;
 END
 END vccdgt_1p0.gds1546
 PIN vccdgt_1p0.gds1547
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.282 27.1435 51.338 27.3435 ;
 END
 END vccdgt_1p0.gds1547
 PIN vccdgt_1p0.gds1548
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.702 26.973 51.758 27.173 ;
 END
 END vccdgt_1p0.gds1548
 PIN vccdgt_1p0.gds1549
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.034 27.163 58.074 27.363 ;
 END
 END vccdgt_1p0.gds1549
 PIN vccdgt_1p0.gds1550
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.762 27.074 57.802 27.274 ;
 END
 END vccdgt_1p0.gds1550
 PIN vccdgt_1p0.gds1551
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.498 27.3135 64.554 27.5135 ;
 END
 END vccdgt_1p0.gds1551
 PIN vccdgt_1p0.gds1552
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.658 27.454 64.714 27.654 ;
 END
 END vccdgt_1p0.gds1552
 PIN vccdgt_1p0.gds1553
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.318 27.119 64.394 27.319 ;
 END
 END vccdgt_1p0.gds1553
 PIN vccdgt_1p0.gds1554
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.834 27.3475 63.874 27.5475 ;
 END
 END vccdgt_1p0.gds1554
 PIN vccdgt_1p0.gds1555
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.158 27.694 65.234 27.894 ;
 END
 END vccdgt_1p0.gds1555
 PIN vccdgt_1p0.gds1556
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.558 27.142 63.618 27.342 ;
 END
 END vccdgt_1p0.gds1556
 PIN vccdgt_1p0.gds1557
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 65.156 27.86 65.212 28.06 ;
 RECT 65.156 26.6 65.212 26.8 ;
 END
 END vccdgt_1p0.gds1557
 PIN vccdgt_1p0.gds1558
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 27.226 67.726 27.426 ;
 END
 END vccdgt_1p0.gds1558
 PIN vccdgt_1p0.gds1559
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 25.966 67.726 26.166 ;
 END
 END vccdgt_1p0.gds1559
 PIN vccdgt_1p0.gds1560
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 28.486 67.726 28.686 ;
 END
 END vccdgt_1p0.gds1560
 PIN vccdgt_1p0.gds1561
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.678 26.9215 65.734 27.1215 ;
 END
 END vccdgt_1p0.gds1561
 PIN vccdgt_1p0.gds1562
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.022 27.5515 67.082 27.7515 ;
 END
 END vccdgt_1p0.gds1562
 PIN vccdgt_1p0.gds1563
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.342 27.5515 66.382 27.7515 ;
 END
 END vccdgt_1p0.gds1563
 PIN vccdgt_1p0.gds1564
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.994 27.9435 68.05 28.1435 ;
 END
 END vccdgt_1p0.gds1564
 PIN vccdgt_1p0.gds1565
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.83 27.6025 67.89 27.8025 ;
 END
 END vccdgt_1p0.gds1565
 PIN vccdgt_1p0.gds1566
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.174 27.936 68.23 28.136 ;
 END
 END vccdgt_1p0.gds1566
 PIN vccdgt_1p0.gds1567
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.494 27.142 68.57 27.342 ;
 END
 END vccdgt_1p0.gds1567
 PIN vccdgt_1p0.gds1568
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.47 27.498 66.51 27.698 ;
 END
 END vccdgt_1p0.gds1568
 PIN vccdgt_1p0.gds1569
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.922 27.036 65.962 27.236 ;
 END
 END vccdgt_1p0.gds1569
 PIN vccdgt_1p0.gds1570
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.338 27.694 65.394 27.894 ;
 END
 END vccdgt_1p0.gds1570
 PIN vccdgt_1p0.gds1571
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.27 27.142 69.33 27.342 ;
 END
 END vccdgt_1p0.gds1571
 PIN vccdgt_1p0.gds1572
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.014 27.984 69.054 28.184 ;
 END
 END vccdgt_1p0.gds1572
 PIN vccdgt_1p0.gds1573
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.334 27.1435 68.39 27.3435 ;
 END
 END vccdgt_1p0.gds1573
 PIN vccdgt_1p0.gds1574
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.114 27.8215 66.154 28.0215 ;
 END
 END vccdgt_1p0.gds1574
 PIN vccdgt_1p0.gds1575
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.754 26.973 68.81 27.173 ;
 END
 END vccdgt_1p0.gds1575
 PIN vccdgt_1p0.gds1576
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.678 27.079 66.738 27.279 ;
 END
 END vccdgt_1p0.gds1576
 PIN vccdgt_1p0.gds1577
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.186 27.709 67.232 27.909 ;
 END
 END vccdgt_1p0.gds1577
 PIN vccdgt_1p0.gds1578
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 65.912 25.457 65.968 25.657 ;
 RECT 67.088 25.52 67.144 25.72 ;
 RECT 65.912 26.717 65.968 26.917 ;
 RECT 67.088 26.78 67.144 26.98 ;
 RECT 65.912 27.977 65.968 28.177 ;
 RECT 67.088 28.04 67.144 28.24 ;
 RECT 66.08 27.544 66.136 27.744 ;
 RECT 66.92 27.62 66.976 27.82 ;
 RECT 66.668 27.872 66.724 28.072 ;
 RECT 66.416 27.959 66.472 28.159 ;
 RECT 65.744 27.977 65.8 28.177 ;
 RECT 67.256 27.977 67.312 28.177 ;
 RECT 65.576 27.964 65.632 28.164 ;
 RECT 66.08 26.284 66.136 26.484 ;
 RECT 66.92 26.36 66.976 26.56 ;
 RECT 66.668 26.612 66.724 26.812 ;
 RECT 66.416 26.699 66.472 26.899 ;
 RECT 65.744 26.717 65.8 26.917 ;
 RECT 67.256 26.717 67.312 26.917 ;
 RECT 65.576 26.704 65.632 26.904 ;
 RECT 65.744 25.457 65.8 25.657 ;
 RECT 67.256 25.457 67.312 25.657 ;
 END
 END vccdgt_1p0.gds1578
END c73p1rfshdxrom2048x16hb4img100_APACHECELL

END LIBRARY
