//=======================================================================
//
// pvr_hqm.vs
//
//
// This module will house the Platfrom Voltage Regulator Module for your
// DUT.  It is to be updated with every voltage domain that is tracked
// and interacted with in your DUT simulations.
//
// Author: <That is you!>
// Date:   <Everyone loves a paper trail>
//
// 
//=======================================================================


//
// Main PVR module for top-level instantiation
//
module pvr_hqm (

  // Inputs
  input real   vcccfn_real,                     // This is the voltage value driven by RTL or TB

  // Outputs
  output logic vcccfn,                          // 0/1 indication to TB/Ascot if Power is on
  output real  vcccfn_on_thresh_out,            // ON  Voltage threshold for driver reference
  output real  vcccfn_ret_thresh_out            // RET Voltage threshold for driver reference

);

// Don't lint the instrumentation code
`ifndef LINT_ON

  ////////////////////////////////////////////////
  //Autogenerated using voltage_instantiation.pl 
  ////////////////////////////////////////////////
  real DOMAIN_VCCCFN_ON_VOLTAGE = 0.65;
  real DOMAIN_VCCCFN_RETENTION_VOLTAGE = 0.30;
  //
  //
  real vcccfn_on_threshold; 
  real vcccfn_ret_threshold; 
  //
  //
  // Threshold initial assignments.  This is done in case fuses or other injections
  // want to run-time override the thresholds.  An example is if a FUSE is used to
  // define the threshold and it is necessary for the Reset Driver to override this
  // value based on that fuse.
  initial begin:PVR_CONST_VOLTAGE
    vcccfn_on_threshold     = DOMAIN_VCCCFN_ON_VOLTAGE; 
    vcccfn_ret_threshold    = DOMAIN_VCCCFN_RETENTION_VOLTAGE; 
  end:PVR_CONST_VOLTAGE

  assign vcccfn_on_thresh_out        = vcccfn_on_threshold;
  assign vcccfn_ret_thresh_out       = vcccfn_ret_threshold;

  //
  //VCCCFN Voltage instantiation
  // - Output:    VCCCFN
  // - INstances:    System
  //
  logic vcccfn_is_retention;
  pvr_voltage_domain #("vcccfn") volt_dom_vcccfn (
    .vcc_out(vcccfn),
    .vcc_retention(vcccfn_is_retention),
    .vcc_in_real(vcccfn_real),
    .vcc_on_voltage(vcccfn_on_threshold),
    .vcc_retention_voltage(vcccfn_ret_threshold),
    .power_enable_in(1)
  );

`endif // LINT_ON

endmodule   // pvr


