// File output was printed on: Wednesday, March 20, 2013 9:00:22 AM
// Chassis TAP Tool version: 0.6.1.2
//----------------------------------------------------------------------
parameter NUMBER_OF_HIER  = 5;
parameter NUMBER_OF_STAPS = 30;
parameter NUMBER_OF_TERTIARY_PORTS = 2;
