interface sbr_par_intf();

logic[15:0] sbr_parity_err_in;
logic       sbr_parity_err_out;
logic[15:0] sbr_port_parity_err;

endinterface
