VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf132b224e1r1w0cbbehcaa4acw
  CLASS BLOCK ;
  FOREIGN arf132b224e1r1w0cbbehcaa4acw ;
  ORIGIN 0 0 ;
  SIZE 79.2 BY 29.76 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.784 16.68 38.828 17.88 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.784 14.76 38.828 15.96 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.86 16.68 39.904 17.88 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.112 16.68 40.156 17.88 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.284 16.68 40.328 17.88 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.872 16.68 38.916 17.88 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.044 16.68 39.088 17.88 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.296 16.68 39.34 17.88 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.472 16.68 39.516 17.88 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.772 16.68 39.816 17.88 ;
    END
  END rdaddrp0[7]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.96 16.68 39.004 17.88 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.212 16.68 39.256 17.88 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.384 16.68 39.428 17.88 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.684 16.68 39.728 17.88 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.112 14.76 40.156 15.96 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.284 14.76 40.328 15.96 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.872 14.76 38.916 15.96 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.044 14.76 39.088 15.96 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.296 14.76 39.34 15.96 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.472 14.76 39.516 15.96 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.772 14.76 39.816 15.96 ;
    END
  END wraddrp0[6]
  PIN wraddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.944 14.76 39.988 15.96 ;
    END
  END wraddrp0[7]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.96 14.76 39.004 15.96 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.212 14.76 39.256 15.96 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.344 0.24 18.388 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 22.56 22.328 23.76 ;
    END
  END wrdatap0[100]
  PIN wrdatap0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 22.56 22.416 23.76 ;
    END
  END wrdatap0[101]
  PIN wrdatap0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.444 22.56 62.488 23.76 ;
    END
  END wrdatap0[102]
  PIN wrdatap0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.528 22.56 62.572 23.76 ;
    END
  END wrdatap0[103]
  PIN wrdatap0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 23.28 18.728 24.48 ;
    END
  END wrdatap0[104]
  PIN wrdatap0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 23.28 18.816 24.48 ;
    END
  END wrdatap0[105]
  PIN wrdatap0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.012 23.28 59.056 24.48 ;
    END
  END wrdatap0[106]
  PIN wrdatap0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.184 23.28 59.228 24.48 ;
    END
  END wrdatap0[107]
  PIN wrdatap0[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 24 20.272 25.2 ;
    END
  END wrdatap0[108]
  PIN wrdatap0[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 24 20.356 25.2 ;
    END
  END wrdatap0[109]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.984 1.68 61.028 2.88 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.384 24 60.428 25.2 ;
    END
  END wrdatap0[110]
  PIN wrdatap0[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.472 24 60.516 25.2 ;
    END
  END wrdatap0[111]
  PIN wrdatap0[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.212 24.72 21.256 25.92 ;
    END
  END wrdatap0[112]
  PIN wrdatap0[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 24.72 21.428 25.92 ;
    END
  END wrdatap0[113]
  PIN wrdatap0[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 24.72 61.416 25.92 ;
    END
  END wrdatap0[114]
  PIN wrdatap0[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.544 24.72 61.588 25.92 ;
    END
  END wrdatap0[115]
  PIN wrdatap0[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 25.44 22.328 26.64 ;
    END
  END wrdatap0[116]
  PIN wrdatap0[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 25.44 22.416 26.64 ;
    END
  END wrdatap0[117]
  PIN wrdatap0[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.444 25.44 62.488 26.64 ;
    END
  END wrdatap0[118]
  PIN wrdatap0[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.528 25.44 62.572 26.64 ;
    END
  END wrdatap0[119]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.072 1.68 61.116 2.88 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 26.16 18.728 27.36 ;
    END
  END wrdatap0[120]
  PIN wrdatap0[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 26.16 18.816 27.36 ;
    END
  END wrdatap0[121]
  PIN wrdatap0[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.012 26.16 59.056 27.36 ;
    END
  END wrdatap0[122]
  PIN wrdatap0[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.184 26.16 59.228 27.36 ;
    END
  END wrdatap0[123]
  PIN wrdatap0[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 26.88 20.272 28.08 ;
    END
  END wrdatap0[124]
  PIN wrdatap0[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 26.88 20.356 28.08 ;
    END
  END wrdatap0[125]
  PIN wrdatap0[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.384 26.88 60.428 28.08 ;
    END
  END wrdatap0[126]
  PIN wrdatap0[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.472 26.88 60.516 28.08 ;
    END
  END wrdatap0[127]
  PIN wrdatap0[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.212 27.6 21.256 28.8 ;
    END
  END wrdatap0[128]
  PIN wrdatap0[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 27.6 21.428 28.8 ;
    END
  END wrdatap0[129]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.944 2.4 21.988 3.6 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 27.6 61.416 28.8 ;
    END
  END wrdatap0[130]
  PIN wrdatap0[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.544 27.6 61.588 28.8 ;
    END
  END wrdatap0[131]
  PIN wrdatap0[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 28.32 22.328 29.52 ;
    END
  END wrdatap0[132]
  PIN wrdatap0[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 28.32 22.416 29.52 ;
    END
  END wrdatap0[133]
  PIN wrdatap0[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.444 28.32 62.488 29.52 ;
    END
  END wrdatap0[134]
  PIN wrdatap0[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.528 28.32 62.572 29.52 ;
    END
  END wrdatap0[135]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 2.4 22.072 3.6 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.972 2.4 62.016 3.6 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.184 2.4 62.228 3.6 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 3.12 22.972 4.32 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 3.12 18.472 4.32 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.372 3.12 58.416 4.32 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.584 3.12 58.628 4.32 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 0.24 18.472 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 3.84 19.716 5.04 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 3.84 19.928 5.04 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.912 3.84 59.956 5.04 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.084 3.84 60.128 5.04 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 4.56 20.916 5.76 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.044 4.56 21.088 5.76 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.984 4.56 61.028 5.76 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.072 4.56 61.116 5.76 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.944 5.28 21.988 6.48 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 5.28 22.072 6.48 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.372 0.24 58.416 1.44 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.972 5.28 62.016 6.48 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.184 5.28 62.228 6.48 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 6 22.972 7.2 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 6 18.472 7.2 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.372 6 58.416 7.2 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.584 6 58.628 7.2 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 6.72 19.716 7.92 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 6.72 19.928 7.92 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.912 6.72 59.956 7.92 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.084 6.72 60.128 7.92 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.584 0.24 58.628 1.44 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 7.44 20.916 8.64 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.044 7.44 21.088 8.64 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.984 7.44 61.028 8.64 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.072 7.44 61.116 8.64 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.944 8.16 21.988 9.36 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 8.16 22.072 9.36 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.972 8.16 62.016 9.36 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.184 8.16 62.228 9.36 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 8.88 22.972 10.08 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 8.88 18.472 10.08 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 0.96 19.928 2.16 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.372 8.88 58.416 10.08 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.584 8.88 58.628 10.08 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 9.6 19.716 10.8 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 9.6 19.928 10.8 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.912 9.6 59.956 10.8 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.084 9.6 60.128 10.8 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 10.32 20.916 11.52 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.044 10.32 21.088 11.52 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.984 10.32 61.028 11.52 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.072 10.32 61.116 11.52 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 0.96 20.016 2.16 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.944 11.04 21.988 12.24 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 11.04 22.072 12.24 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.972 11.04 62.016 12.24 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.184 11.04 62.228 12.24 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 11.76 22.972 12.96 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 11.76 18.472 12.96 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.372 11.76 58.416 12.96 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.584 11.76 58.628 12.96 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 12.48 19.716 13.68 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 12.48 19.928 13.68 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.912 0.96 59.956 2.16 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.912 12.48 59.956 13.68 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.084 12.48 60.128 13.68 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 13.2 20.916 14.4 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.044 13.2 21.088 14.4 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.984 13.2 61.028 14.4 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.072 13.2 61.116 14.4 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 18.24 19.716 19.44 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 18.24 19.928 19.44 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.828 18.24 59.872 19.44 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.912 18.24 59.956 19.44 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.084 0.96 60.128 2.16 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.212 18.96 21.256 20.16 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 18.96 21.428 20.16 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 18.96 61.416 20.16 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.544 18.96 61.588 20.16 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 19.68 22.328 20.88 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 19.68 22.416 20.88 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.444 19.68 62.488 20.88 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.528 19.68 62.572 20.88 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 20.4 18.728 21.6 ;
    END
  END wrdatap0[88]
  PIN wrdatap0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 20.4 18.816 21.6 ;
    END
  END wrdatap0[89]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 1.68 20.916 2.88 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.012 20.4 59.056 21.6 ;
    END
  END wrdatap0[90]
  PIN wrdatap0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.184 20.4 59.228 21.6 ;
    END
  END wrdatap0[91]
  PIN wrdatap0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 21.12 20.272 22.32 ;
    END
  END wrdatap0[92]
  PIN wrdatap0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 21.12 20.356 22.32 ;
    END
  END wrdatap0[93]
  PIN wrdatap0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.384 21.12 60.428 22.32 ;
    END
  END wrdatap0[94]
  PIN wrdatap0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.472 21.12 60.516 22.32 ;
    END
  END wrdatap0[95]
  PIN wrdatap0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.212 21.84 21.256 23.04 ;
    END
  END wrdatap0[96]
  PIN wrdatap0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 21.84 21.428 23.04 ;
    END
  END wrdatap0[97]
  PIN wrdatap0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 21.84 61.416 23.04 ;
    END
  END wrdatap0[98]
  PIN wrdatap0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.544 21.84 61.588 23.04 ;
    END
  END wrdatap0[99]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.044 1.68 21.088 2.88 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.684 14.76 39.728 15.96 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.86 14.76 39.904 15.96 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.384 14.76 39.428 15.96 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 0.24 18.556 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 22.56 22.628 23.76 ;
    END
  END rddatap0[100]
  PIN rddatap0[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 22.56 22.716 23.76 ;
    END
  END rddatap0[101]
  PIN rddatap0[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.028 22.56 58.072 23.76 ;
    END
  END rddatap0[102]
  PIN rddatap0[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.112 22.56 58.156 23.76 ;
    END
  END rddatap0[103]
  PIN rddatap0[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 23.28 19.028 24.48 ;
    END
  END rddatap0[104]
  PIN rddatap0[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 23.28 19.116 24.48 ;
    END
  END rddatap0[105]
  PIN rddatap0[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.272 23.28 59.316 24.48 ;
    END
  END rddatap0[106]
  PIN rddatap0[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.484 23.28 59.528 24.48 ;
    END
  END rddatap0[107]
  PIN rddatap0[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 24 20.528 25.2 ;
    END
  END rddatap0[108]
  PIN rddatap0[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 24 20.616 25.2 ;
    END
  END rddatap0[109]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.284 1.68 61.328 2.88 ;
    END
  END rddatap0[10]
  PIN rddatap0[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.644 24 60.688 25.2 ;
    END
  END rddatap0[110]
  PIN rddatap0[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.728 24 60.772 25.2 ;
    END
  END rddatap0[111]
  PIN rddatap0[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 24.72 21.516 25.92 ;
    END
  END rddatap0[112]
  PIN rddatap0[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 24.72 21.728 25.92 ;
    END
  END rddatap0[113]
  PIN rddatap0[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.628 24.72 61.672 25.92 ;
    END
  END rddatap0[114]
  PIN rddatap0[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.712 24.72 61.756 25.92 ;
    END
  END rddatap0[115]
  PIN rddatap0[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 25.44 22.628 26.64 ;
    END
  END rddatap0[116]
  PIN rddatap0[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 25.44 22.716 26.64 ;
    END
  END rddatap0[117]
  PIN rddatap0[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.028 25.44 58.072 26.64 ;
    END
  END rddatap0[118]
  PIN rddatap0[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.112 25.44 58.156 26.64 ;
    END
  END rddatap0[119]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 1.68 61.416 2.88 ;
    END
  END rddatap0[11]
  PIN rddatap0[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 26.16 19.028 27.36 ;
    END
  END rddatap0[120]
  PIN rddatap0[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 26.16 19.116 27.36 ;
    END
  END rddatap0[121]
  PIN rddatap0[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.272 26.16 59.316 27.36 ;
    END
  END rddatap0[122]
  PIN rddatap0[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.484 26.16 59.528 27.36 ;
    END
  END rddatap0[123]
  PIN rddatap0[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 26.88 20.528 28.08 ;
    END
  END rddatap0[124]
  PIN rddatap0[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 26.88 20.616 28.08 ;
    END
  END rddatap0[125]
  PIN rddatap0[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.644 26.88 60.688 28.08 ;
    END
  END rddatap0[126]
  PIN rddatap0[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.728 26.88 60.772 28.08 ;
    END
  END rddatap0[127]
  PIN rddatap0[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 27.6 21.516 28.8 ;
    END
  END rddatap0[128]
  PIN rddatap0[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 27.6 21.728 28.8 ;
    END
  END rddatap0[129]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.112 2.4 22.156 3.6 ;
    END
  END rddatap0[12]
  PIN rddatap0[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.628 27.6 61.672 28.8 ;
    END
  END rddatap0[130]
  PIN rddatap0[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.712 27.6 61.756 28.8 ;
    END
  END rddatap0[131]
  PIN rddatap0[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 28.32 22.628 29.52 ;
    END
  END rddatap0[132]
  PIN rddatap0[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 28.32 22.716 29.52 ;
    END
  END rddatap0[133]
  PIN rddatap0[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.028 28.32 58.072 29.52 ;
    END
  END rddatap0[134]
  PIN rddatap0[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.112 28.32 58.156 29.52 ;
    END
  END rddatap0[135]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 2.4 22.328 3.6 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.272 2.4 62.316 3.6 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.444 2.4 62.488 3.6 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 3.12 18.556 4.32 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 3.12 18.728 4.32 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.672 3.12 58.716 4.32 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.844 3.12 58.888 4.32 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 0.24 18.728 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 3.84 20.016 5.04 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.144 3.84 20.188 5.04 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.172 3.84 60.216 5.04 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.384 3.84 60.428 5.04 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 4.56 21.172 5.76 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.212 4.56 21.256 5.76 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.284 4.56 61.328 5.76 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 4.56 61.416 5.76 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.112 5.28 22.156 6.48 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 5.28 22.328 6.48 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.672 0.24 58.716 1.44 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.272 5.28 62.316 6.48 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.444 5.28 62.488 6.48 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 6 18.556 7.2 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 6 18.728 7.2 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.672 6 58.716 7.2 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.844 6 58.888 7.2 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 6.72 20.016 7.92 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.144 6.72 20.188 7.92 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.172 6.72 60.216 7.92 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.384 6.72 60.428 7.92 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.844 0.24 58.888 1.44 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 7.44 21.172 8.64 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.212 7.44 21.256 8.64 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.284 7.44 61.328 8.64 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 7.44 61.416 8.64 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.112 8.16 22.156 9.36 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 8.16 22.328 9.36 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.272 8.16 62.316 9.36 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.444 8.16 62.488 9.36 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 8.88 18.556 10.08 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 8.88 18.728 10.08 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.144 0.96 20.188 2.16 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.672 8.88 58.716 10.08 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.844 8.88 58.888 10.08 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 9.6 20.016 10.8 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.144 9.6 20.188 10.8 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.172 9.6 60.216 10.8 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.384 9.6 60.428 10.8 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 10.32 21.172 11.52 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.212 10.32 21.256 11.52 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.284 10.32 61.328 11.52 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 10.32 61.416 11.52 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 0.96 20.272 2.16 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.112 11.04 22.156 12.24 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 11.04 22.328 12.24 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.272 11.04 62.316 12.24 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.444 11.04 62.488 12.24 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 11.76 18.556 12.96 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 11.76 18.728 12.96 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.672 11.76 58.716 12.96 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.844 11.76 58.888 12.96 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 12.48 20.016 13.68 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.144 12.48 20.188 13.68 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.172 0.96 60.216 2.16 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.172 12.48 60.216 13.68 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.384 12.48 60.428 13.68 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 13.2 21.172 14.4 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.212 13.2 21.256 14.4 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.284 13.2 61.328 14.4 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 13.2 61.416 14.4 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 18.24 20.016 19.44 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.144 18.24 20.188 19.44 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.084 18.24 60.128 19.44 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.172 18.24 60.216 19.44 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.384 0.96 60.428 2.16 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 18.96 21.516 20.16 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 18.96 21.728 20.16 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.628 18.96 61.672 20.16 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.712 18.96 61.756 20.16 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 19.68 22.628 20.88 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 19.68 22.716 20.88 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.028 19.68 58.072 20.88 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 58.112 19.68 58.156 20.88 ;
    END
  END rddatap0[87]
  PIN rddatap0[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 20.4 19.028 21.6 ;
    END
  END rddatap0[88]
  PIN rddatap0[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 20.4 19.116 21.6 ;
    END
  END rddatap0[89]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 1.68 21.172 2.88 ;
    END
  END rddatap0[8]
  PIN rddatap0[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.272 20.4 59.316 21.6 ;
    END
  END rddatap0[90]
  PIN rddatap0[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 59.484 20.4 59.528 21.6 ;
    END
  END rddatap0[91]
  PIN rddatap0[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 21.12 20.528 22.32 ;
    END
  END rddatap0[92]
  PIN rddatap0[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 21.12 20.616 22.32 ;
    END
  END rddatap0[93]
  PIN rddatap0[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.644 21.12 60.688 22.32 ;
    END
  END rddatap0[94]
  PIN rddatap0[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 60.728 21.12 60.772 22.32 ;
    END
  END rddatap0[95]
  PIN rddatap0[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 21.84 21.516 23.04 ;
    END
  END rddatap0[96]
  PIN rddatap0[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 21.84 21.728 23.04 ;
    END
  END rddatap0[97]
  PIN rddatap0[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.628 21.84 61.672 23.04 ;
    END
  END rddatap0[98]
  PIN rddatap0[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.712 21.84 61.756 23.04 ;
    END
  END rddatap0[99]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.212 1.68 21.256 2.88 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 29.7 ;
        RECT 2.662 0.06 2.738 29.7 ;
        RECT 4.462 0.06 4.538 29.7 ;
        RECT 6.262 0.06 6.338 29.7 ;
        RECT 8.062 0.06 8.138 29.7 ;
        RECT 9.862 0.06 9.938 29.7 ;
        RECT 11.662 0.06 11.738 29.7 ;
        RECT 13.462 0.06 13.538 29.7 ;
        RECT 15.262 0.06 15.338 29.7 ;
        RECT 17.062 0.06 17.138 29.7 ;
        RECT 18.862 0.06 18.938 29.7 ;
        RECT 20.662 0.06 20.738 29.7 ;
        RECT 22.462 0.06 22.538 29.7 ;
        RECT 24.262 0.06 24.338 29.7 ;
        RECT 26.062 0.06 26.138 29.7 ;
        RECT 27.862 0.06 27.938 29.7 ;
        RECT 29.662 0.06 29.738 29.7 ;
        RECT 31.462 0.06 31.538 29.7 ;
        RECT 33.262 0.06 33.338 29.7 ;
        RECT 35.062 0.06 35.138 29.7 ;
        RECT 36.862 0.06 36.938 29.7 ;
        RECT 38.662 0.06 38.738 29.7 ;
        RECT 40.462 0.06 40.538 29.7 ;
        RECT 42.262 0.06 42.338 29.7 ;
        RECT 44.062 0.06 44.138 29.7 ;
        RECT 45.862 0.06 45.938 29.7 ;
        RECT 47.662 0.06 47.738 29.7 ;
        RECT 49.462 0.06 49.538 29.7 ;
        RECT 51.262 0.06 51.338 29.7 ;
        RECT 53.062 0.06 53.138 29.7 ;
        RECT 54.862 0.06 54.938 29.7 ;
        RECT 56.662 0.06 56.738 29.7 ;
        RECT 58.462 0.06 58.538 29.7 ;
        RECT 60.262 0.06 60.338 29.7 ;
        RECT 62.062 0.06 62.138 29.7 ;
        RECT 63.862 0.06 63.938 29.7 ;
        RECT 65.662 0.06 65.738 29.7 ;
        RECT 67.462 0.06 67.538 29.7 ;
        RECT 69.262 0.06 69.338 29.7 ;
        RECT 71.062 0.06 71.138 29.7 ;
        RECT 72.862 0.06 72.938 29.7 ;
        RECT 74.662 0.06 74.738 29.7 ;
        RECT 76.462 0.06 76.538 29.7 ;
        RECT 78.262 0.06 78.338 29.7 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 29.7 ;
        RECT 3.562 0.06 3.638 29.7 ;
        RECT 5.362 0.06 5.438 29.7 ;
        RECT 7.162 0.06 7.238 29.7 ;
        RECT 8.962 0.06 9.038 29.7 ;
        RECT 10.762 0.06 10.838 29.7 ;
        RECT 12.562 0.06 12.638 29.7 ;
        RECT 14.362 0.06 14.438 29.7 ;
        RECT 16.162 0.06 16.238 29.7 ;
        RECT 17.962 0.06 18.038 29.7 ;
        RECT 19.762 0.06 19.838 29.7 ;
        RECT 21.562 0.06 21.638 29.7 ;
        RECT 23.362 0.06 23.438 29.7 ;
        RECT 25.162 0.06 25.238 29.7 ;
        RECT 26.962 0.06 27.038 29.7 ;
        RECT 28.762 0.06 28.838 29.7 ;
        RECT 30.562 0.06 30.638 29.7 ;
        RECT 32.362 0.06 32.438 29.7 ;
        RECT 34.162 0.06 34.238 29.7 ;
        RECT 35.962 0.06 36.038 29.7 ;
        RECT 37.762 0.06 37.838 29.7 ;
        RECT 39.562 0.06 39.638 29.7 ;
        RECT 41.362 0.06 41.438 29.7 ;
        RECT 43.162 0.06 43.238 29.7 ;
        RECT 44.962 0.06 45.038 29.7 ;
        RECT 46.762 0.06 46.838 29.7 ;
        RECT 48.562 0.06 48.638 29.7 ;
        RECT 50.362 0.06 50.438 29.7 ;
        RECT 52.162 0.06 52.238 29.7 ;
        RECT 53.962 0.06 54.038 29.7 ;
        RECT 55.762 0.06 55.838 29.7 ;
        RECT 57.562 0.06 57.638 29.7 ;
        RECT 59.362 0.06 59.438 29.7 ;
        RECT 61.162 0.06 61.238 29.7 ;
        RECT 62.962 0.06 63.038 29.7 ;
        RECT 64.762 0.06 64.838 29.7 ;
        RECT 66.562 0.06 66.638 29.7 ;
        RECT 68.362 0.06 68.438 29.7 ;
        RECT 70.162 0.06 70.238 29.7 ;
        RECT 71.962 0.06 72.038 29.7 ;
        RECT 73.762 0.06 73.838 29.7 ;
        RECT 75.562 0.06 75.638 29.7 ;
        RECT 77.362 0.06 77.438 29.7 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 79.216 29.774 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 79.22 29.78 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 79.2705 29.798 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 79.235 29.83 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 79.27 29.798 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 79.259 29.85 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 79.29 29.822 ;
    LAYER m7 SPACING 0 ;
      RECT 78.338 29.82 79.24 29.88 ;
      RECT 78.338 -0.06 79.292 29.82 ;
      RECT 78.338 -0.12 79.24 -0.06 ;
      RECT 77.438 -0.12 78.262 29.88 ;
      RECT 76.538 -0.12 77.362 29.88 ;
      RECT 75.638 -0.12 76.462 29.88 ;
      RECT 74.738 -0.12 75.562 29.88 ;
      RECT 73.838 -0.12 74.662 29.88 ;
      RECT 72.938 -0.12 73.762 29.88 ;
      RECT 72.038 -0.12 72.862 29.88 ;
      RECT 71.138 -0.12 71.962 29.88 ;
      RECT 70.238 -0.12 71.062 29.88 ;
      RECT 69.338 -0.12 70.162 29.88 ;
      RECT 68.438 -0.12 69.262 29.88 ;
      RECT 67.538 -0.12 68.362 29.88 ;
      RECT 66.638 -0.12 67.462 29.88 ;
      RECT 65.738 -0.12 66.562 29.88 ;
      RECT 64.838 -0.12 65.662 29.88 ;
      RECT 63.938 -0.12 64.762 29.88 ;
      RECT 63.038 -0.12 63.862 29.88 ;
      RECT 62.138 29.52 62.962 29.88 ;
      RECT 62.138 28.32 62.444 29.52 ;
      RECT 62.488 28.32 62.528 29.52 ;
      RECT 62.572 28.32 62.962 29.52 ;
      RECT 62.138 26.64 62.962 28.32 ;
      RECT 62.138 25.44 62.444 26.64 ;
      RECT 62.488 25.44 62.528 26.64 ;
      RECT 62.572 25.44 62.962 26.64 ;
      RECT 62.138 23.76 62.962 25.44 ;
      RECT 62.138 22.56 62.444 23.76 ;
      RECT 62.488 22.56 62.528 23.76 ;
      RECT 62.572 22.56 62.962 23.76 ;
      RECT 62.138 20.88 62.962 22.56 ;
      RECT 62.138 19.68 62.444 20.88 ;
      RECT 62.488 19.68 62.528 20.88 ;
      RECT 62.572 19.68 62.962 20.88 ;
      RECT 62.138 12.24 62.962 19.68 ;
      RECT 62.138 11.04 62.184 12.24 ;
      RECT 62.228 11.04 62.272 12.24 ;
      RECT 62.316 11.04 62.444 12.24 ;
      RECT 62.488 11.04 62.962 12.24 ;
      RECT 62.138 9.36 62.962 11.04 ;
      RECT 62.138 8.16 62.184 9.36 ;
      RECT 62.228 8.16 62.272 9.36 ;
      RECT 62.316 8.16 62.444 9.36 ;
      RECT 62.488 8.16 62.962 9.36 ;
      RECT 62.138 6.48 62.962 8.16 ;
      RECT 62.138 5.28 62.184 6.48 ;
      RECT 62.228 5.28 62.272 6.48 ;
      RECT 62.316 5.28 62.444 6.48 ;
      RECT 62.488 5.28 62.962 6.48 ;
      RECT 62.138 3.6 62.962 5.28 ;
      RECT 62.138 2.4 62.184 3.6 ;
      RECT 62.228 2.4 62.272 3.6 ;
      RECT 62.316 2.4 62.444 3.6 ;
      RECT 62.488 2.4 62.962 3.6 ;
      RECT 62.138 -0.12 62.962 2.4 ;
      RECT 61.238 28.8 62.062 29.88 ;
      RECT 61.238 27.6 61.372 28.8 ;
      RECT 61.416 27.6 61.544 28.8 ;
      RECT 61.588 27.6 61.628 28.8 ;
      RECT 61.672 27.6 61.712 28.8 ;
      RECT 61.756 27.6 62.062 28.8 ;
      RECT 61.238 25.92 62.062 27.6 ;
      RECT 61.238 24.72 61.372 25.92 ;
      RECT 61.416 24.72 61.544 25.92 ;
      RECT 61.588 24.72 61.628 25.92 ;
      RECT 61.672 24.72 61.712 25.92 ;
      RECT 61.756 24.72 62.062 25.92 ;
      RECT 61.238 23.04 62.062 24.72 ;
      RECT 61.238 21.84 61.372 23.04 ;
      RECT 61.416 21.84 61.544 23.04 ;
      RECT 61.588 21.84 61.628 23.04 ;
      RECT 61.672 21.84 61.712 23.04 ;
      RECT 61.756 21.84 62.062 23.04 ;
      RECT 61.238 20.16 62.062 21.84 ;
      RECT 61.238 18.96 61.372 20.16 ;
      RECT 61.416 18.96 61.544 20.16 ;
      RECT 61.588 18.96 61.628 20.16 ;
      RECT 61.672 18.96 61.712 20.16 ;
      RECT 61.756 18.96 62.062 20.16 ;
      RECT 61.238 14.4 62.062 18.96 ;
      RECT 61.238 13.2 61.284 14.4 ;
      RECT 61.328 13.2 61.372 14.4 ;
      RECT 61.416 13.2 62.062 14.4 ;
      RECT 61.238 12.24 62.062 13.2 ;
      RECT 61.238 11.52 61.972 12.24 ;
      RECT 62.016 11.04 62.062 12.24 ;
      RECT 61.416 11.04 61.972 11.52 ;
      RECT 61.238 10.32 61.284 11.52 ;
      RECT 61.328 10.32 61.372 11.52 ;
      RECT 61.416 10.32 62.062 11.04 ;
      RECT 61.238 9.36 62.062 10.32 ;
      RECT 61.238 8.64 61.972 9.36 ;
      RECT 62.016 8.16 62.062 9.36 ;
      RECT 61.416 8.16 61.972 8.64 ;
      RECT 61.238 7.44 61.284 8.64 ;
      RECT 61.328 7.44 61.372 8.64 ;
      RECT 61.416 7.44 62.062 8.16 ;
      RECT 61.238 6.48 62.062 7.44 ;
      RECT 61.238 5.76 61.972 6.48 ;
      RECT 62.016 5.28 62.062 6.48 ;
      RECT 61.416 5.28 61.972 5.76 ;
      RECT 61.238 4.56 61.284 5.76 ;
      RECT 61.328 4.56 61.372 5.76 ;
      RECT 61.416 4.56 62.062 5.28 ;
      RECT 61.238 3.6 62.062 4.56 ;
      RECT 61.238 2.88 61.972 3.6 ;
      RECT 62.016 2.4 62.062 3.6 ;
      RECT 61.416 2.4 61.972 2.88 ;
      RECT 61.238 1.68 61.284 2.88 ;
      RECT 61.328 1.68 61.372 2.88 ;
      RECT 61.416 1.68 62.062 2.4 ;
      RECT 61.238 -0.12 62.062 1.68 ;
      RECT 60.338 28.08 61.162 29.88 ;
      RECT 60.338 26.88 60.384 28.08 ;
      RECT 60.428 26.88 60.472 28.08 ;
      RECT 60.516 26.88 60.644 28.08 ;
      RECT 60.688 26.88 60.728 28.08 ;
      RECT 60.772 26.88 61.162 28.08 ;
      RECT 60.338 25.2 61.162 26.88 ;
      RECT 60.338 24 60.384 25.2 ;
      RECT 60.428 24 60.472 25.2 ;
      RECT 60.516 24 60.644 25.2 ;
      RECT 60.688 24 60.728 25.2 ;
      RECT 60.772 24 61.162 25.2 ;
      RECT 60.338 22.32 61.162 24 ;
      RECT 60.338 21.12 60.384 22.32 ;
      RECT 60.428 21.12 60.472 22.32 ;
      RECT 60.516 21.12 60.644 22.32 ;
      RECT 60.688 21.12 60.728 22.32 ;
      RECT 60.772 21.12 61.162 22.32 ;
      RECT 60.338 14.4 61.162 21.12 ;
      RECT 60.338 13.68 60.984 14.4 ;
      RECT 61.028 13.2 61.072 14.4 ;
      RECT 61.116 13.2 61.162 14.4 ;
      RECT 60.428 13.2 60.984 13.68 ;
      RECT 60.338 12.48 60.384 13.68 ;
      RECT 60.428 12.48 61.162 13.2 ;
      RECT 60.338 11.52 61.162 12.48 ;
      RECT 60.338 10.8 60.984 11.52 ;
      RECT 61.028 10.32 61.072 11.52 ;
      RECT 61.116 10.32 61.162 11.52 ;
      RECT 60.428 10.32 60.984 10.8 ;
      RECT 60.338 9.6 60.384 10.8 ;
      RECT 60.428 9.6 61.162 10.32 ;
      RECT 60.338 8.64 61.162 9.6 ;
      RECT 60.338 7.92 60.984 8.64 ;
      RECT 61.028 7.44 61.072 8.64 ;
      RECT 61.116 7.44 61.162 8.64 ;
      RECT 60.428 7.44 60.984 7.92 ;
      RECT 60.338 6.72 60.384 7.92 ;
      RECT 60.428 6.72 61.162 7.44 ;
      RECT 60.338 5.76 61.162 6.72 ;
      RECT 60.338 5.04 60.984 5.76 ;
      RECT 61.028 4.56 61.072 5.76 ;
      RECT 61.116 4.56 61.162 5.76 ;
      RECT 60.428 4.56 60.984 5.04 ;
      RECT 60.338 3.84 60.384 5.04 ;
      RECT 60.428 3.84 61.162 4.56 ;
      RECT 60.338 2.88 61.162 3.84 ;
      RECT 60.338 2.16 60.984 2.88 ;
      RECT 61.028 1.68 61.072 2.88 ;
      RECT 61.116 1.68 61.162 2.88 ;
      RECT 60.428 1.68 60.984 2.16 ;
      RECT 60.338 0.96 60.384 2.16 ;
      RECT 60.428 0.96 61.162 1.68 ;
      RECT 60.338 -0.12 61.162 0.96 ;
      RECT 59.438 27.36 60.262 29.88 ;
      RECT 59.438 26.16 59.484 27.36 ;
      RECT 59.528 26.16 60.262 27.36 ;
      RECT 59.438 24.48 60.262 26.16 ;
      RECT 59.438 23.28 59.484 24.48 ;
      RECT 59.528 23.28 60.262 24.48 ;
      RECT 59.438 21.6 60.262 23.28 ;
      RECT 59.438 20.4 59.484 21.6 ;
      RECT 59.528 20.4 60.262 21.6 ;
      RECT 59.438 19.44 60.262 20.4 ;
      RECT 59.438 18.24 59.828 19.44 ;
      RECT 59.872 18.24 59.912 19.44 ;
      RECT 59.956 18.24 60.084 19.44 ;
      RECT 60.128 18.24 60.172 19.44 ;
      RECT 60.216 18.24 60.262 19.44 ;
      RECT 59.438 13.68 60.262 18.24 ;
      RECT 59.438 12.48 59.912 13.68 ;
      RECT 59.956 12.48 60.084 13.68 ;
      RECT 60.128 12.48 60.172 13.68 ;
      RECT 60.216 12.48 60.262 13.68 ;
      RECT 59.438 10.8 60.262 12.48 ;
      RECT 59.438 9.6 59.912 10.8 ;
      RECT 59.956 9.6 60.084 10.8 ;
      RECT 60.128 9.6 60.172 10.8 ;
      RECT 60.216 9.6 60.262 10.8 ;
      RECT 59.438 7.92 60.262 9.6 ;
      RECT 59.438 6.72 59.912 7.92 ;
      RECT 59.956 6.72 60.084 7.92 ;
      RECT 60.128 6.72 60.172 7.92 ;
      RECT 60.216 6.72 60.262 7.92 ;
      RECT 59.438 5.04 60.262 6.72 ;
      RECT 59.438 3.84 59.912 5.04 ;
      RECT 59.956 3.84 60.084 5.04 ;
      RECT 60.128 3.84 60.172 5.04 ;
      RECT 60.216 3.84 60.262 5.04 ;
      RECT 59.438 2.16 60.262 3.84 ;
      RECT 59.438 0.96 59.912 2.16 ;
      RECT 59.956 0.96 60.084 2.16 ;
      RECT 60.128 0.96 60.172 2.16 ;
      RECT 60.216 0.96 60.262 2.16 ;
      RECT 59.438 -0.12 60.262 0.96 ;
      RECT 58.538 27.36 59.362 29.88 ;
      RECT 58.538 26.16 59.012 27.36 ;
      RECT 59.056 26.16 59.184 27.36 ;
      RECT 59.228 26.16 59.272 27.36 ;
      RECT 59.316 26.16 59.362 27.36 ;
      RECT 58.538 24.48 59.362 26.16 ;
      RECT 58.538 23.28 59.012 24.48 ;
      RECT 59.056 23.28 59.184 24.48 ;
      RECT 59.228 23.28 59.272 24.48 ;
      RECT 59.316 23.28 59.362 24.48 ;
      RECT 58.538 21.6 59.362 23.28 ;
      RECT 58.538 20.4 59.012 21.6 ;
      RECT 59.056 20.4 59.184 21.6 ;
      RECT 59.228 20.4 59.272 21.6 ;
      RECT 59.316 20.4 59.362 21.6 ;
      RECT 58.538 12.96 59.362 20.4 ;
      RECT 58.538 11.76 58.584 12.96 ;
      RECT 58.628 11.76 58.672 12.96 ;
      RECT 58.716 11.76 58.844 12.96 ;
      RECT 58.888 11.76 59.362 12.96 ;
      RECT 58.538 10.08 59.362 11.76 ;
      RECT 58.538 8.88 58.584 10.08 ;
      RECT 58.628 8.88 58.672 10.08 ;
      RECT 58.716 8.88 58.844 10.08 ;
      RECT 58.888 8.88 59.362 10.08 ;
      RECT 58.538 7.2 59.362 8.88 ;
      RECT 58.538 6 58.584 7.2 ;
      RECT 58.628 6 58.672 7.2 ;
      RECT 58.716 6 58.844 7.2 ;
      RECT 58.888 6 59.362 7.2 ;
      RECT 58.538 4.32 59.362 6 ;
      RECT 58.538 3.12 58.584 4.32 ;
      RECT 58.628 3.12 58.672 4.32 ;
      RECT 58.716 3.12 58.844 4.32 ;
      RECT 58.888 3.12 59.362 4.32 ;
      RECT 58.538 1.44 59.362 3.12 ;
      RECT 58.538 0.24 58.584 1.44 ;
      RECT 58.628 0.24 58.672 1.44 ;
      RECT 58.716 0.24 58.844 1.44 ;
      RECT 58.888 0.24 59.362 1.44 ;
      RECT 58.538 -0.12 59.362 0.24 ;
      RECT 57.638 29.52 58.462 29.88 ;
      RECT 57.638 28.32 58.028 29.52 ;
      RECT 58.072 28.32 58.112 29.52 ;
      RECT 58.156 28.32 58.462 29.52 ;
      RECT 57.638 26.64 58.462 28.32 ;
      RECT 57.638 25.44 58.028 26.64 ;
      RECT 58.072 25.44 58.112 26.64 ;
      RECT 58.156 25.44 58.462 26.64 ;
      RECT 57.638 23.76 58.462 25.44 ;
      RECT 57.638 22.56 58.028 23.76 ;
      RECT 58.072 22.56 58.112 23.76 ;
      RECT 58.156 22.56 58.462 23.76 ;
      RECT 57.638 20.88 58.462 22.56 ;
      RECT 57.638 19.68 58.028 20.88 ;
      RECT 58.072 19.68 58.112 20.88 ;
      RECT 58.156 19.68 58.462 20.88 ;
      RECT 57.638 12.96 58.462 19.68 ;
      RECT 57.638 11.76 58.372 12.96 ;
      RECT 58.416 11.76 58.462 12.96 ;
      RECT 57.638 10.08 58.462 11.76 ;
      RECT 57.638 8.88 58.372 10.08 ;
      RECT 58.416 8.88 58.462 10.08 ;
      RECT 57.638 7.2 58.462 8.88 ;
      RECT 57.638 6 58.372 7.2 ;
      RECT 58.416 6 58.462 7.2 ;
      RECT 57.638 4.32 58.462 6 ;
      RECT 57.638 3.12 58.372 4.32 ;
      RECT 58.416 3.12 58.462 4.32 ;
      RECT 57.638 1.44 58.462 3.12 ;
      RECT 57.638 0.24 58.372 1.44 ;
      RECT 58.416 0.24 58.462 1.44 ;
      RECT 57.638 -0.12 58.462 0.24 ;
      RECT 56.738 -0.12 57.562 29.88 ;
      RECT 55.838 -0.12 56.662 29.88 ;
      RECT 54.938 -0.12 55.762 29.88 ;
      RECT 54.038 -0.12 54.862 29.88 ;
      RECT 53.138 -0.12 53.962 29.88 ;
      RECT 52.238 -0.12 53.062 29.88 ;
      RECT 51.338 -0.12 52.162 29.88 ;
      RECT 50.438 -0.12 51.262 29.88 ;
      RECT 49.538 -0.12 50.362 29.88 ;
      RECT 48.638 -0.12 49.462 29.88 ;
      RECT 47.738 -0.12 48.562 29.88 ;
      RECT 46.838 -0.12 47.662 29.88 ;
      RECT 45.938 -0.12 46.762 29.88 ;
      RECT 45.038 -0.12 45.862 29.88 ;
      RECT 44.138 -0.12 44.962 29.88 ;
      RECT 43.238 -0.12 44.062 29.88 ;
      RECT 42.338 -0.12 43.162 29.88 ;
      RECT 41.438 -0.12 42.262 29.88 ;
      RECT 40.538 -0.12 41.362 29.88 ;
      RECT 39.638 17.88 40.462 29.88 ;
      RECT 39.638 16.68 39.684 17.88 ;
      RECT 39.728 16.68 39.772 17.88 ;
      RECT 39.816 16.68 39.86 17.88 ;
      RECT 39.904 16.68 40.112 17.88 ;
      RECT 40.156 16.68 40.284 17.88 ;
      RECT 40.328 16.68 40.462 17.88 ;
      RECT 39.638 15.96 40.462 16.68 ;
      RECT 39.638 14.76 39.684 15.96 ;
      RECT 39.728 14.76 39.772 15.96 ;
      RECT 39.816 14.76 39.86 15.96 ;
      RECT 39.904 14.76 39.944 15.96 ;
      RECT 39.988 14.76 40.112 15.96 ;
      RECT 40.156 14.76 40.284 15.96 ;
      RECT 40.328 14.76 40.462 15.96 ;
      RECT 39.638 -0.12 40.462 14.76 ;
      RECT 38.738 17.88 39.562 29.88 ;
      RECT 38.738 16.68 38.784 17.88 ;
      RECT 38.828 16.68 38.872 17.88 ;
      RECT 38.916 16.68 38.96 17.88 ;
      RECT 39.004 16.68 39.044 17.88 ;
      RECT 39.088 16.68 39.212 17.88 ;
      RECT 39.256 16.68 39.296 17.88 ;
      RECT 39.34 16.68 39.384 17.88 ;
      RECT 39.428 16.68 39.472 17.88 ;
      RECT 39.516 16.68 39.562 17.88 ;
      RECT 38.738 15.96 39.562 16.68 ;
      RECT 38.738 14.76 38.784 15.96 ;
      RECT 38.828 14.76 38.872 15.96 ;
      RECT 38.916 14.76 38.96 15.96 ;
      RECT 39.004 14.76 39.044 15.96 ;
      RECT 39.088 14.76 39.212 15.96 ;
      RECT 39.256 14.76 39.296 15.96 ;
      RECT 39.34 14.76 39.384 15.96 ;
      RECT 39.428 14.76 39.472 15.96 ;
      RECT 39.516 14.76 39.562 15.96 ;
      RECT 38.738 -0.12 39.562 14.76 ;
      RECT 37.838 -0.12 38.662 29.88 ;
      RECT 36.938 -0.12 37.762 29.88 ;
      RECT 36.038 -0.12 36.862 29.88 ;
      RECT 35.138 -0.12 35.962 29.88 ;
      RECT 34.238 -0.12 35.062 29.88 ;
      RECT 33.338 -0.12 34.162 29.88 ;
      RECT 32.438 -0.12 33.262 29.88 ;
      RECT 31.538 -0.12 32.362 29.88 ;
      RECT 30.638 -0.12 31.462 29.88 ;
      RECT 29.738 -0.12 30.562 29.88 ;
      RECT 28.838 -0.12 29.662 29.88 ;
      RECT 27.938 -0.12 28.762 29.88 ;
      RECT 27.038 -0.12 27.862 29.88 ;
      RECT 26.138 -0.12 26.962 29.88 ;
      RECT 25.238 -0.12 26.062 29.88 ;
      RECT 24.338 -0.12 25.162 29.88 ;
      RECT 23.438 -0.12 24.262 29.88 ;
      RECT 22.538 29.52 23.362 29.88 ;
      RECT 22.538 28.32 22.584 29.52 ;
      RECT 22.628 28.32 22.672 29.52 ;
      RECT 22.716 28.32 23.362 29.52 ;
      RECT 22.538 26.64 23.362 28.32 ;
      RECT 22.538 25.44 22.584 26.64 ;
      RECT 22.628 25.44 22.672 26.64 ;
      RECT 22.716 25.44 23.362 26.64 ;
      RECT 22.538 23.76 23.362 25.44 ;
      RECT 22.538 22.56 22.584 23.76 ;
      RECT 22.628 22.56 22.672 23.76 ;
      RECT 22.716 22.56 23.362 23.76 ;
      RECT 22.538 20.88 23.362 22.56 ;
      RECT 22.538 19.68 22.584 20.88 ;
      RECT 22.628 19.68 22.672 20.88 ;
      RECT 22.716 19.68 23.362 20.88 ;
      RECT 22.538 12.96 23.362 19.68 ;
      RECT 22.538 11.76 22.928 12.96 ;
      RECT 22.972 11.76 23.362 12.96 ;
      RECT 22.538 10.08 23.362 11.76 ;
      RECT 22.538 8.88 22.928 10.08 ;
      RECT 22.972 8.88 23.362 10.08 ;
      RECT 22.538 7.2 23.362 8.88 ;
      RECT 22.538 6 22.928 7.2 ;
      RECT 22.972 6 23.362 7.2 ;
      RECT 22.538 4.32 23.362 6 ;
      RECT 22.538 3.12 22.928 4.32 ;
      RECT 22.972 3.12 23.362 4.32 ;
      RECT 22.538 -0.12 23.362 3.12 ;
      RECT 21.638 29.52 22.462 29.88 ;
      RECT 21.638 28.8 22.284 29.52 ;
      RECT 22.328 28.32 22.372 29.52 ;
      RECT 22.416 28.32 22.462 29.52 ;
      RECT 21.728 28.32 22.284 28.8 ;
      RECT 21.638 27.6 21.684 28.8 ;
      RECT 21.728 27.6 22.462 28.32 ;
      RECT 21.638 26.64 22.462 27.6 ;
      RECT 21.638 25.92 22.284 26.64 ;
      RECT 22.328 25.44 22.372 26.64 ;
      RECT 22.416 25.44 22.462 26.64 ;
      RECT 21.728 25.44 22.284 25.92 ;
      RECT 21.638 24.72 21.684 25.92 ;
      RECT 21.728 24.72 22.462 25.44 ;
      RECT 21.638 23.76 22.462 24.72 ;
      RECT 21.638 23.04 22.284 23.76 ;
      RECT 22.328 22.56 22.372 23.76 ;
      RECT 22.416 22.56 22.462 23.76 ;
      RECT 21.728 22.56 22.284 23.04 ;
      RECT 21.638 21.84 21.684 23.04 ;
      RECT 21.728 21.84 22.462 22.56 ;
      RECT 21.638 20.88 22.462 21.84 ;
      RECT 21.638 20.16 22.284 20.88 ;
      RECT 22.328 19.68 22.372 20.88 ;
      RECT 22.416 19.68 22.462 20.88 ;
      RECT 21.728 19.68 22.284 20.16 ;
      RECT 21.638 18.96 21.684 20.16 ;
      RECT 21.728 18.96 22.462 19.68 ;
      RECT 21.638 12.24 22.462 18.96 ;
      RECT 21.638 11.04 21.944 12.24 ;
      RECT 21.988 11.04 22.028 12.24 ;
      RECT 22.072 11.04 22.112 12.24 ;
      RECT 22.156 11.04 22.284 12.24 ;
      RECT 22.328 11.04 22.462 12.24 ;
      RECT 21.638 9.36 22.462 11.04 ;
      RECT 21.638 8.16 21.944 9.36 ;
      RECT 21.988 8.16 22.028 9.36 ;
      RECT 22.072 8.16 22.112 9.36 ;
      RECT 22.156 8.16 22.284 9.36 ;
      RECT 22.328 8.16 22.462 9.36 ;
      RECT 21.638 6.48 22.462 8.16 ;
      RECT 21.638 5.28 21.944 6.48 ;
      RECT 21.988 5.28 22.028 6.48 ;
      RECT 22.072 5.28 22.112 6.48 ;
      RECT 22.156 5.28 22.284 6.48 ;
      RECT 22.328 5.28 22.462 6.48 ;
      RECT 21.638 3.6 22.462 5.28 ;
      RECT 21.638 2.4 21.944 3.6 ;
      RECT 21.988 2.4 22.028 3.6 ;
      RECT 22.072 2.4 22.112 3.6 ;
      RECT 22.156 2.4 22.284 3.6 ;
      RECT 22.328 2.4 22.462 3.6 ;
      RECT 21.638 -0.12 22.462 2.4 ;
      RECT 20.738 28.8 21.562 29.88 ;
      RECT 20.738 27.6 21.212 28.8 ;
      RECT 21.256 27.6 21.384 28.8 ;
      RECT 21.428 27.6 21.472 28.8 ;
      RECT 21.516 27.6 21.562 28.8 ;
      RECT 20.738 25.92 21.562 27.6 ;
      RECT 20.738 24.72 21.212 25.92 ;
      RECT 21.256 24.72 21.384 25.92 ;
      RECT 21.428 24.72 21.472 25.92 ;
      RECT 21.516 24.72 21.562 25.92 ;
      RECT 20.738 23.04 21.562 24.72 ;
      RECT 20.738 21.84 21.212 23.04 ;
      RECT 21.256 21.84 21.384 23.04 ;
      RECT 21.428 21.84 21.472 23.04 ;
      RECT 21.516 21.84 21.562 23.04 ;
      RECT 20.738 20.16 21.562 21.84 ;
      RECT 20.738 18.96 21.212 20.16 ;
      RECT 21.256 18.96 21.384 20.16 ;
      RECT 21.428 18.96 21.472 20.16 ;
      RECT 21.516 18.96 21.562 20.16 ;
      RECT 20.738 14.4 21.562 18.96 ;
      RECT 20.738 13.2 20.872 14.4 ;
      RECT 20.916 13.2 21.044 14.4 ;
      RECT 21.088 13.2 21.128 14.4 ;
      RECT 21.172 13.2 21.212 14.4 ;
      RECT 21.256 13.2 21.562 14.4 ;
      RECT 20.738 11.52 21.562 13.2 ;
      RECT 20.738 10.32 20.872 11.52 ;
      RECT 20.916 10.32 21.044 11.52 ;
      RECT 21.088 10.32 21.128 11.52 ;
      RECT 21.172 10.32 21.212 11.52 ;
      RECT 21.256 10.32 21.562 11.52 ;
      RECT 20.738 8.64 21.562 10.32 ;
      RECT 20.738 7.44 20.872 8.64 ;
      RECT 20.916 7.44 21.044 8.64 ;
      RECT 21.088 7.44 21.128 8.64 ;
      RECT 21.172 7.44 21.212 8.64 ;
      RECT 21.256 7.44 21.562 8.64 ;
      RECT 20.738 5.76 21.562 7.44 ;
      RECT 20.738 4.56 20.872 5.76 ;
      RECT 20.916 4.56 21.044 5.76 ;
      RECT 21.088 4.56 21.128 5.76 ;
      RECT 21.172 4.56 21.212 5.76 ;
      RECT 21.256 4.56 21.562 5.76 ;
      RECT 20.738 2.88 21.562 4.56 ;
      RECT 20.738 1.68 20.872 2.88 ;
      RECT 20.916 1.68 21.044 2.88 ;
      RECT 21.088 1.68 21.128 2.88 ;
      RECT 21.172 1.68 21.212 2.88 ;
      RECT 21.256 1.68 21.562 2.88 ;
      RECT 20.738 -0.12 21.562 1.68 ;
      RECT 19.838 28.08 20.662 29.88 ;
      RECT 19.838 26.88 20.228 28.08 ;
      RECT 20.272 26.88 20.312 28.08 ;
      RECT 20.356 26.88 20.484 28.08 ;
      RECT 20.528 26.88 20.572 28.08 ;
      RECT 20.616 26.88 20.662 28.08 ;
      RECT 19.838 25.2 20.662 26.88 ;
      RECT 19.838 24 20.228 25.2 ;
      RECT 20.272 24 20.312 25.2 ;
      RECT 20.356 24 20.484 25.2 ;
      RECT 20.528 24 20.572 25.2 ;
      RECT 20.616 24 20.662 25.2 ;
      RECT 19.838 22.32 20.662 24 ;
      RECT 19.838 21.12 20.228 22.32 ;
      RECT 20.272 21.12 20.312 22.32 ;
      RECT 20.356 21.12 20.484 22.32 ;
      RECT 20.528 21.12 20.572 22.32 ;
      RECT 20.616 21.12 20.662 22.32 ;
      RECT 19.838 19.44 20.662 21.12 ;
      RECT 19.838 18.24 19.884 19.44 ;
      RECT 19.928 18.24 19.972 19.44 ;
      RECT 20.016 18.24 20.144 19.44 ;
      RECT 20.188 18.24 20.662 19.44 ;
      RECT 19.838 13.68 20.662 18.24 ;
      RECT 19.838 12.48 19.884 13.68 ;
      RECT 19.928 12.48 19.972 13.68 ;
      RECT 20.016 12.48 20.144 13.68 ;
      RECT 20.188 12.48 20.662 13.68 ;
      RECT 19.838 10.8 20.662 12.48 ;
      RECT 19.838 9.6 19.884 10.8 ;
      RECT 19.928 9.6 19.972 10.8 ;
      RECT 20.016 9.6 20.144 10.8 ;
      RECT 20.188 9.6 20.662 10.8 ;
      RECT 19.838 7.92 20.662 9.6 ;
      RECT 19.838 6.72 19.884 7.92 ;
      RECT 19.928 6.72 19.972 7.92 ;
      RECT 20.016 6.72 20.144 7.92 ;
      RECT 20.188 6.72 20.662 7.92 ;
      RECT 19.838 5.04 20.662 6.72 ;
      RECT 19.838 3.84 19.884 5.04 ;
      RECT 19.928 3.84 19.972 5.04 ;
      RECT 20.016 3.84 20.144 5.04 ;
      RECT 20.188 3.84 20.662 5.04 ;
      RECT 19.838 2.16 20.662 3.84 ;
      RECT 19.838 0.96 19.884 2.16 ;
      RECT 19.928 0.96 19.972 2.16 ;
      RECT 20.016 0.96 20.144 2.16 ;
      RECT 20.188 0.96 20.228 2.16 ;
      RECT 20.272 0.96 20.662 2.16 ;
      RECT 19.838 -0.12 20.662 0.96 ;
      RECT 18.938 27.36 19.762 29.88 ;
      RECT 18.938 26.16 18.984 27.36 ;
      RECT 19.028 26.16 19.072 27.36 ;
      RECT 19.116 26.16 19.762 27.36 ;
      RECT 18.938 24.48 19.762 26.16 ;
      RECT 18.938 23.28 18.984 24.48 ;
      RECT 19.028 23.28 19.072 24.48 ;
      RECT 19.116 23.28 19.762 24.48 ;
      RECT 18.938 21.6 19.762 23.28 ;
      RECT 18.938 20.4 18.984 21.6 ;
      RECT 19.028 20.4 19.072 21.6 ;
      RECT 19.116 20.4 19.762 21.6 ;
      RECT 18.938 19.44 19.762 20.4 ;
      RECT 18.938 18.24 19.672 19.44 ;
      RECT 19.716 18.24 19.762 19.44 ;
      RECT 18.938 13.68 19.762 18.24 ;
      RECT 18.938 12.48 19.672 13.68 ;
      RECT 19.716 12.48 19.762 13.68 ;
      RECT 18.938 10.8 19.762 12.48 ;
      RECT 18.938 9.6 19.672 10.8 ;
      RECT 19.716 9.6 19.762 10.8 ;
      RECT 18.938 7.92 19.762 9.6 ;
      RECT 18.938 6.72 19.672 7.92 ;
      RECT 19.716 6.72 19.762 7.92 ;
      RECT 18.938 5.04 19.762 6.72 ;
      RECT 18.938 3.84 19.672 5.04 ;
      RECT 19.716 3.84 19.762 5.04 ;
      RECT 18.938 -0.12 19.762 3.84 ;
      RECT 18.038 27.36 18.862 29.88 ;
      RECT 18.038 26.16 18.684 27.36 ;
      RECT 18.728 26.16 18.772 27.36 ;
      RECT 18.816 26.16 18.862 27.36 ;
      RECT 18.038 24.48 18.862 26.16 ;
      RECT 18.038 23.28 18.684 24.48 ;
      RECT 18.728 23.28 18.772 24.48 ;
      RECT 18.816 23.28 18.862 24.48 ;
      RECT 18.038 21.6 18.862 23.28 ;
      RECT 18.038 20.4 18.684 21.6 ;
      RECT 18.728 20.4 18.772 21.6 ;
      RECT 18.816 20.4 18.862 21.6 ;
      RECT 18.038 12.96 18.862 20.4 ;
      RECT 18.038 11.76 18.428 12.96 ;
      RECT 18.472 11.76 18.512 12.96 ;
      RECT 18.556 11.76 18.684 12.96 ;
      RECT 18.728 11.76 18.862 12.96 ;
      RECT 18.038 10.08 18.862 11.76 ;
      RECT 18.038 8.88 18.428 10.08 ;
      RECT 18.472 8.88 18.512 10.08 ;
      RECT 18.556 8.88 18.684 10.08 ;
      RECT 18.728 8.88 18.862 10.08 ;
      RECT 18.038 7.2 18.862 8.88 ;
      RECT 18.038 6 18.428 7.2 ;
      RECT 18.472 6 18.512 7.2 ;
      RECT 18.556 6 18.684 7.2 ;
      RECT 18.728 6 18.862 7.2 ;
      RECT 18.038 4.32 18.862 6 ;
      RECT 18.038 3.12 18.428 4.32 ;
      RECT 18.472 3.12 18.512 4.32 ;
      RECT 18.556 3.12 18.684 4.32 ;
      RECT 18.728 3.12 18.862 4.32 ;
      RECT 18.038 1.44 18.862 3.12 ;
      RECT 18.038 0.24 18.344 1.44 ;
      RECT 18.388 0.24 18.428 1.44 ;
      RECT 18.472 0.24 18.512 1.44 ;
      RECT 18.556 0.24 18.684 1.44 ;
      RECT 18.728 0.24 18.862 1.44 ;
      RECT 18.038 -0.12 18.862 0.24 ;
      RECT 17.138 -0.12 17.962 29.88 ;
      RECT 16.238 -0.12 17.062 29.88 ;
      RECT 15.338 -0.12 16.162 29.88 ;
      RECT 14.438 -0.12 15.262 29.88 ;
      RECT 13.538 -0.12 14.362 29.88 ;
      RECT 12.638 -0.12 13.462 29.88 ;
      RECT 11.738 -0.12 12.562 29.88 ;
      RECT 10.838 -0.12 11.662 29.88 ;
      RECT 9.938 -0.12 10.762 29.88 ;
      RECT 9.038 -0.12 9.862 29.88 ;
      RECT 8.138 -0.12 8.962 29.88 ;
      RECT 7.238 -0.12 8.062 29.88 ;
      RECT 6.338 -0.12 7.162 29.88 ;
      RECT 5.438 -0.12 6.262 29.88 ;
      RECT 4.538 -0.12 5.362 29.88 ;
      RECT 3.638 -0.12 4.462 29.88 ;
      RECT 2.738 -0.12 3.562 29.88 ;
      RECT 1.838 -0.12 2.662 29.88 ;
      RECT 0.938 -0.12 1.762 29.88 ;
      RECT -0.04 29.82 0.862 29.88 ;
      RECT -0.092 -0.06 0.862 29.82 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 78.458 0 79.12 29.76 ;
      RECT 77.558 0 78.142 29.76 ;
      RECT 76.658 0 77.242 29.76 ;
      RECT 75.758 0 76.342 29.76 ;
      RECT 74.858 0 75.442 29.76 ;
      RECT 73.958 0 74.542 29.76 ;
      RECT 73.058 0 73.642 29.76 ;
      RECT 72.158 0 72.742 29.76 ;
      RECT 71.258 0 71.842 29.76 ;
      RECT 70.358 0 70.942 29.76 ;
      RECT 69.458 0 70.042 29.76 ;
      RECT 68.558 0 69.142 29.76 ;
      RECT 67.658 0 68.242 29.76 ;
      RECT 66.758 0 67.342 29.76 ;
      RECT 65.858 0 66.442 29.76 ;
      RECT 64.958 0 65.542 29.76 ;
      RECT 64.058 0 64.642 29.76 ;
      RECT 63.158 0 63.742 29.76 ;
      RECT 62.258 29.64 62.842 29.76 ;
      RECT 62.258 28.2 62.324 29.64 ;
      RECT 62.692 28.2 62.842 29.64 ;
      RECT 62.258 26.76 62.842 28.2 ;
      RECT 62.258 25.32 62.324 26.76 ;
      RECT 62.692 25.32 62.842 26.76 ;
      RECT 62.258 23.88 62.842 25.32 ;
      RECT 62.258 22.44 62.324 23.88 ;
      RECT 62.692 22.44 62.842 23.88 ;
      RECT 62.258 21 62.842 22.44 ;
      RECT 62.258 19.56 62.324 21 ;
      RECT 62.692 19.56 62.842 21 ;
      RECT 62.258 12.36 62.842 19.56 ;
      RECT 62.608 10.92 62.842 12.36 ;
      RECT 62.258 9.48 62.842 10.92 ;
      RECT 62.608 8.04 62.842 9.48 ;
      RECT 62.258 6.6 62.842 8.04 ;
      RECT 62.608 5.16 62.842 6.6 ;
      RECT 62.258 3.72 62.842 5.16 ;
      RECT 62.608 2.28 62.842 3.72 ;
      RECT 62.258 0 62.842 2.28 ;
      RECT 61.358 28.92 61.942 29.76 ;
      RECT 61.876 27.48 61.942 28.92 ;
      RECT 61.358 26.04 61.942 27.48 ;
      RECT 61.876 24.6 61.942 26.04 ;
      RECT 61.358 23.16 61.942 24.6 ;
      RECT 61.876 21.72 61.942 23.16 ;
      RECT 61.358 20.28 61.942 21.72 ;
      RECT 61.876 18.84 61.942 20.28 ;
      RECT 61.358 14.52 61.942 18.84 ;
      RECT 61.536 13.08 61.942 14.52 ;
      RECT 61.358 12.36 61.942 13.08 ;
      RECT 61.358 11.64 61.852 12.36 ;
      RECT 61.536 10.92 61.852 11.64 ;
      RECT 61.536 10.2 61.942 10.92 ;
      RECT 61.358 9.48 61.942 10.2 ;
      RECT 61.358 8.76 61.852 9.48 ;
      RECT 61.536 8.04 61.852 8.76 ;
      RECT 61.536 7.32 61.942 8.04 ;
      RECT 61.358 6.6 61.942 7.32 ;
      RECT 61.358 5.88 61.852 6.6 ;
      RECT 61.536 5.16 61.852 5.88 ;
      RECT 61.536 4.44 61.942 5.16 ;
      RECT 61.358 3.72 61.942 4.44 ;
      RECT 61.358 3 61.852 3.72 ;
      RECT 61.536 2.28 61.852 3 ;
      RECT 61.536 1.56 61.942 2.28 ;
      RECT 61.358 0 61.942 1.56 ;
      RECT 60.458 28.2 61.042 29.76 ;
      RECT 60.892 26.76 61.042 28.2 ;
      RECT 60.458 25.32 61.042 26.76 ;
      RECT 60.892 23.88 61.042 25.32 ;
      RECT 60.458 22.44 61.042 23.88 ;
      RECT 60.892 21 61.042 22.44 ;
      RECT 60.458 14.52 61.042 21 ;
      RECT 60.458 13.8 60.864 14.52 ;
      RECT 60.548 13.08 60.864 13.8 ;
      RECT 60.548 12.36 61.042 13.08 ;
      RECT 60.458 11.64 61.042 12.36 ;
      RECT 60.458 10.92 60.864 11.64 ;
      RECT 60.548 10.2 60.864 10.92 ;
      RECT 60.548 9.48 61.042 10.2 ;
      RECT 60.458 8.76 61.042 9.48 ;
      RECT 60.458 8.04 60.864 8.76 ;
      RECT 60.548 7.32 60.864 8.04 ;
      RECT 60.548 6.6 61.042 7.32 ;
      RECT 60.458 5.88 61.042 6.6 ;
      RECT 60.458 5.16 60.864 5.88 ;
      RECT 60.548 4.44 60.864 5.16 ;
      RECT 60.548 3.72 61.042 4.44 ;
      RECT 60.458 3 61.042 3.72 ;
      RECT 60.458 2.28 60.864 3 ;
      RECT 60.548 1.56 60.864 2.28 ;
      RECT 60.548 0.84 61.042 1.56 ;
      RECT 60.458 0 61.042 0.84 ;
      RECT 59.558 27.48 60.142 29.76 ;
      RECT 59.648 26.04 60.142 27.48 ;
      RECT 59.558 24.6 60.142 26.04 ;
      RECT 59.648 23.16 60.142 24.6 ;
      RECT 59.558 21.72 60.142 23.16 ;
      RECT 59.648 20.28 60.142 21.72 ;
      RECT 59.558 19.56 60.142 20.28 ;
      RECT 59.558 18.12 59.708 19.56 ;
      RECT 59.558 13.8 60.142 18.12 ;
      RECT 59.558 12.36 59.792 13.8 ;
      RECT 59.558 10.92 60.142 12.36 ;
      RECT 59.558 9.48 59.792 10.92 ;
      RECT 59.558 8.04 60.142 9.48 ;
      RECT 59.558 6.6 59.792 8.04 ;
      RECT 59.558 5.16 60.142 6.6 ;
      RECT 59.558 3.72 59.792 5.16 ;
      RECT 59.558 2.28 60.142 3.72 ;
      RECT 59.558 0.84 59.792 2.28 ;
      RECT 59.558 0 60.142 0.84 ;
      RECT 58.658 27.48 59.242 29.76 ;
      RECT 58.658 26.04 58.892 27.48 ;
      RECT 58.658 24.6 59.242 26.04 ;
      RECT 58.658 23.16 58.892 24.6 ;
      RECT 58.658 21.72 59.242 23.16 ;
      RECT 58.658 20.28 58.892 21.72 ;
      RECT 58.658 13.08 59.242 20.28 ;
      RECT 59.008 11.64 59.242 13.08 ;
      RECT 58.658 10.2 59.242 11.64 ;
      RECT 59.008 8.76 59.242 10.2 ;
      RECT 58.658 7.32 59.242 8.76 ;
      RECT 59.008 5.88 59.242 7.32 ;
      RECT 58.658 4.44 59.242 5.88 ;
      RECT 59.008 3 59.242 4.44 ;
      RECT 58.658 1.56 59.242 3 ;
      RECT 59.008 0.12 59.242 1.56 ;
      RECT 58.658 0 59.242 0.12 ;
      RECT 57.758 29.64 58.342 29.76 ;
      RECT 57.758 28.2 57.908 29.64 ;
      RECT 58.276 28.2 58.342 29.64 ;
      RECT 57.758 26.76 58.342 28.2 ;
      RECT 57.758 25.32 57.908 26.76 ;
      RECT 58.276 25.32 58.342 26.76 ;
      RECT 57.758 23.88 58.342 25.32 ;
      RECT 57.758 22.44 57.908 23.88 ;
      RECT 58.276 22.44 58.342 23.88 ;
      RECT 57.758 21 58.342 22.44 ;
      RECT 57.758 19.56 57.908 21 ;
      RECT 58.276 19.56 58.342 21 ;
      RECT 57.758 13.08 58.342 19.56 ;
      RECT 57.758 11.64 58.252 13.08 ;
      RECT 57.758 10.2 58.342 11.64 ;
      RECT 57.758 8.76 58.252 10.2 ;
      RECT 57.758 7.32 58.342 8.76 ;
      RECT 57.758 5.88 58.252 7.32 ;
      RECT 57.758 4.44 58.342 5.88 ;
      RECT 57.758 3 58.252 4.44 ;
      RECT 57.758 1.56 58.342 3 ;
      RECT 57.758 0.12 58.252 1.56 ;
      RECT 57.758 0 58.342 0.12 ;
      RECT 56.858 0 57.442 29.76 ;
      RECT 55.958 0 56.542 29.76 ;
      RECT 55.058 0 55.642 29.76 ;
      RECT 54.158 0 54.742 29.76 ;
      RECT 53.258 0 53.842 29.76 ;
      RECT 52.358 0 52.942 29.76 ;
      RECT 51.458 0 52.042 29.76 ;
      RECT 50.558 0 51.142 29.76 ;
      RECT 49.658 0 50.242 29.76 ;
      RECT 48.758 0 49.342 29.76 ;
      RECT 47.858 0 48.442 29.76 ;
      RECT 46.958 0 47.542 29.76 ;
      RECT 46.058 0 46.642 29.76 ;
      RECT 45.158 0 45.742 29.76 ;
      RECT 44.258 0 44.842 29.76 ;
      RECT 43.358 0 43.942 29.76 ;
      RECT 42.458 0 43.042 29.76 ;
      RECT 41.558 0 42.142 29.76 ;
      RECT 40.658 0 41.242 29.76 ;
      RECT 39.758 18 40.342 29.76 ;
      RECT 38.858 18 39.442 29.76 ;
      RECT 37.958 0 38.542 29.76 ;
      RECT 37.058 0 37.642 29.76 ;
      RECT 36.158 0 36.742 29.76 ;
      RECT 35.258 0 35.842 29.76 ;
      RECT 34.358 0 34.942 29.76 ;
      RECT 33.458 0 34.042 29.76 ;
      RECT 32.558 0 33.142 29.76 ;
      RECT 31.658 0 32.242 29.76 ;
      RECT 30.758 0 31.342 29.76 ;
      RECT 29.858 0 30.442 29.76 ;
      RECT 28.958 0 29.542 29.76 ;
      RECT 28.058 0 28.642 29.76 ;
      RECT 27.158 0 27.742 29.76 ;
      RECT 26.258 0 26.842 29.76 ;
      RECT 25.358 0 25.942 29.76 ;
      RECT 24.458 0 25.042 29.76 ;
      RECT 23.558 0 24.142 29.76 ;
      RECT 22.658 29.64 23.242 29.76 ;
      RECT 22.836 28.2 23.242 29.64 ;
      RECT 22.658 26.76 23.242 28.2 ;
      RECT 22.836 25.32 23.242 26.76 ;
      RECT 22.658 23.88 23.242 25.32 ;
      RECT 22.836 22.44 23.242 23.88 ;
      RECT 22.658 21 23.242 22.44 ;
      RECT 22.836 19.56 23.242 21 ;
      RECT 22.658 13.08 23.242 19.56 ;
      RECT 22.658 11.64 22.808 13.08 ;
      RECT 23.092 11.64 23.242 13.08 ;
      RECT 22.658 10.2 23.242 11.64 ;
      RECT 22.658 8.76 22.808 10.2 ;
      RECT 23.092 8.76 23.242 10.2 ;
      RECT 22.658 7.32 23.242 8.76 ;
      RECT 22.658 5.88 22.808 7.32 ;
      RECT 23.092 5.88 23.242 7.32 ;
      RECT 22.658 4.44 23.242 5.88 ;
      RECT 22.658 3 22.808 4.44 ;
      RECT 23.092 3 23.242 4.44 ;
      RECT 22.658 0 23.242 3 ;
      RECT 21.758 29.64 22.342 29.76 ;
      RECT 21.758 28.92 22.164 29.64 ;
      RECT 21.848 28.2 22.164 28.92 ;
      RECT 21.848 27.48 22.342 28.2 ;
      RECT 21.758 26.76 22.342 27.48 ;
      RECT 21.758 26.04 22.164 26.76 ;
      RECT 21.848 25.32 22.164 26.04 ;
      RECT 21.848 24.6 22.342 25.32 ;
      RECT 21.758 23.88 22.342 24.6 ;
      RECT 21.758 23.16 22.164 23.88 ;
      RECT 21.848 22.44 22.164 23.16 ;
      RECT 21.848 21.72 22.342 22.44 ;
      RECT 21.758 21 22.342 21.72 ;
      RECT 21.758 20.28 22.164 21 ;
      RECT 21.848 19.56 22.164 20.28 ;
      RECT 21.848 18.84 22.342 19.56 ;
      RECT 21.758 12.36 22.342 18.84 ;
      RECT 21.758 10.92 21.824 12.36 ;
      RECT 21.758 9.48 22.342 10.92 ;
      RECT 21.758 8.04 21.824 9.48 ;
      RECT 21.758 6.6 22.342 8.04 ;
      RECT 21.758 5.16 21.824 6.6 ;
      RECT 21.758 3.72 22.342 5.16 ;
      RECT 21.758 2.28 21.824 3.72 ;
      RECT 21.758 0 22.342 2.28 ;
      RECT 20.858 28.92 21.442 29.76 ;
      RECT 20.858 27.48 21.092 28.92 ;
      RECT 20.858 26.04 21.442 27.48 ;
      RECT 20.858 24.6 21.092 26.04 ;
      RECT 20.858 23.16 21.442 24.6 ;
      RECT 20.858 21.72 21.092 23.16 ;
      RECT 20.858 20.28 21.442 21.72 ;
      RECT 20.858 18.84 21.092 20.28 ;
      RECT 20.858 14.52 21.442 18.84 ;
      RECT 21.376 13.08 21.442 14.52 ;
      RECT 20.858 11.64 21.442 13.08 ;
      RECT 21.376 10.2 21.442 11.64 ;
      RECT 20.858 8.76 21.442 10.2 ;
      RECT 21.376 7.32 21.442 8.76 ;
      RECT 20.858 5.88 21.442 7.32 ;
      RECT 21.376 4.44 21.442 5.88 ;
      RECT 20.858 3 21.442 4.44 ;
      RECT 21.376 1.56 21.442 3 ;
      RECT 20.858 0 21.442 1.56 ;
      RECT 19.958 28.2 20.542 29.76 ;
      RECT 19.958 26.76 20.108 28.2 ;
      RECT 19.958 25.32 20.542 26.76 ;
      RECT 19.958 23.88 20.108 25.32 ;
      RECT 19.958 22.44 20.542 23.88 ;
      RECT 19.958 21 20.108 22.44 ;
      RECT 19.958 19.56 20.542 21 ;
      RECT 20.308 18.12 20.542 19.56 ;
      RECT 19.958 13.8 20.542 18.12 ;
      RECT 20.308 12.36 20.542 13.8 ;
      RECT 19.958 10.92 20.542 12.36 ;
      RECT 20.308 9.48 20.542 10.92 ;
      RECT 19.958 8.04 20.542 9.48 ;
      RECT 20.308 6.6 20.542 8.04 ;
      RECT 19.958 5.16 20.542 6.6 ;
      RECT 20.308 3.72 20.542 5.16 ;
      RECT 19.958 2.28 20.542 3.72 ;
      RECT 20.392 0.84 20.542 2.28 ;
      RECT 19.958 0 20.542 0.84 ;
      RECT 19.058 27.48 19.642 29.76 ;
      RECT 19.236 26.04 19.642 27.48 ;
      RECT 19.058 24.6 19.642 26.04 ;
      RECT 19.236 23.16 19.642 24.6 ;
      RECT 19.058 21.72 19.642 23.16 ;
      RECT 19.236 20.28 19.642 21.72 ;
      RECT 19.058 19.56 19.642 20.28 ;
      RECT 19.058 18.12 19.552 19.56 ;
      RECT 19.058 13.8 19.642 18.12 ;
      RECT 19.058 12.36 19.552 13.8 ;
      RECT 19.058 10.92 19.642 12.36 ;
      RECT 19.058 9.48 19.552 10.92 ;
      RECT 19.058 8.04 19.642 9.48 ;
      RECT 19.058 6.6 19.552 8.04 ;
      RECT 19.058 5.16 19.642 6.6 ;
      RECT 19.058 3.72 19.552 5.16 ;
      RECT 19.058 0 19.642 3.72 ;
      RECT 18.158 27.48 18.742 29.76 ;
      RECT 18.158 26.04 18.564 27.48 ;
      RECT 18.158 24.6 18.742 26.04 ;
      RECT 18.158 23.16 18.564 24.6 ;
      RECT 18.158 21.72 18.742 23.16 ;
      RECT 18.158 20.28 18.564 21.72 ;
      RECT 18.158 13.08 18.742 20.28 ;
      RECT 18.158 11.64 18.308 13.08 ;
      RECT 18.158 10.2 18.742 11.64 ;
      RECT 18.158 8.76 18.308 10.2 ;
      RECT 18.158 7.32 18.742 8.76 ;
      RECT 18.158 5.88 18.308 7.32 ;
      RECT 18.158 4.44 18.742 5.88 ;
      RECT 18.158 3 18.308 4.44 ;
      RECT 18.158 1.56 18.742 3 ;
      RECT 18.158 0.12 18.224 1.56 ;
      RECT 18.158 0 18.742 0.12 ;
      RECT 17.258 0 17.842 29.76 ;
      RECT 16.358 0 16.942 29.76 ;
      RECT 15.458 0 16.042 29.76 ;
      RECT 14.558 0 15.142 29.76 ;
      RECT 13.658 0 14.242 29.76 ;
      RECT 12.758 0 13.342 29.76 ;
      RECT 11.858 0 12.442 29.76 ;
      RECT 10.958 0 11.542 29.76 ;
      RECT 10.058 0 10.642 29.76 ;
      RECT 9.158 0 9.742 29.76 ;
      RECT 8.258 0 8.842 29.76 ;
      RECT 7.358 0 7.942 29.76 ;
      RECT 6.458 0 7.042 29.76 ;
      RECT 5.558 0 6.142 29.76 ;
      RECT 4.658 0 5.242 29.76 ;
      RECT 3.758 0 4.342 29.76 ;
      RECT 2.858 0 3.442 29.76 ;
      RECT 1.958 0 2.542 29.76 ;
      RECT 1.058 0 1.642 29.76 ;
      RECT 0.08 0 0.742 29.76 ;
      RECT 39.758 16.08 40.342 16.56 ;
      RECT 38.858 16.08 39.442 16.56 ;
      RECT 39.758 0 40.342 14.64 ;
      RECT 38.858 0 39.442 14.64 ;
    LAYER m0 ;
      RECT 0 0.002 79.2 29.758 ;
    LAYER m1 ;
      RECT 0 0 79.2 29.76 ;
    LAYER m2 ;
      RECT 0 0.015 79.2 29.745 ;
    LAYER m3 ;
      RECT 0.015 0 79.185 29.76 ;
    LAYER m4 ;
      RECT 0 0.02 79.2 29.74 ;
    LAYER m5 ;
      RECT 0.012 0 79.188 29.76 ;
    LAYER m6 ;
      RECT 0 0.012 79.2 29.748 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf132b224e1r1w0cbbehcaa4acw

END LIBRARY
