// RTL Generated using Collage

module hqm_sip_aon_wrap # (
    // Subsystem Parameters
    parameter HQM_DTF_DATA_WIDTH = 64,
    parameter HQM_DTF_HEADER_WIDTH = 25,
    parameter HQM_DTF_TO_CNT_THRESHOLD = 1000,
    parameter HQM_DVP_USE_LEGACY_TIMESTAMP = 0,
    parameter HQM_DVP_USE_PUSH_SWD = 0,
    parameter HQM_SBE_DATAWIDTH = 8,
    parameter HQM_SBE_NPQUEUEDEPTH = 4,
    parameter HQM_SBE_PARITY_REQUIRED = 1,
    parameter HQM_SBE_PCQUEUEDEPTH = 4,
    parameter HQM_SFI_RX_BCM_EN = 1,
    parameter HQM_SFI_RX_BLOCK_EARLY_VLD_EN = 1,
    parameter HQM_SFI_RX_D = 32,
    parameter HQM_SFI_RX_DATA_AUX_PARITY_EN = 1,
    parameter HQM_SFI_RX_DATA_CRD_GRAN = 4,
    parameter HQM_SFI_RX_DATA_INTERLEAVE = 0,
    parameter HQM_SFI_RX_DATA_LAYER_EN = 1,
    parameter HQM_SFI_RX_DATA_MAX_FC_VC = 1,
    parameter HQM_SFI_RX_DATA_PARITY_EN = 1,
    parameter HQM_SFI_RX_DATA_PASS_HDR = 0,
    parameter HQM_SFI_RX_DS = 1,
    parameter HQM_SFI_RX_ECRC_SUPPORT = 0,
    parameter HQM_SFI_RX_FATAL_EN = 0,
    parameter HQM_SFI_RX_FLIT_MODE_PREFIX_EN = 0,
    parameter HQM_SFI_RX_H = 32,
    parameter HQM_SFI_RX_HDR_DATA_SEP = 1,
    parameter HQM_SFI_RX_HDR_MAX_FC_VC = 1,
    parameter HQM_SFI_RX_HGRAN = 4,
    parameter HQM_SFI_RX_HPARITY = 1,
    parameter HQM_SFI_RX_IDE_SUPPORT = 0,
    parameter HQM_SFI_RX_M = 1,
    parameter HQM_SFI_RX_MAX_CRD_CNT_WIDTH = 12,
    parameter HQM_SFI_RX_MAX_HDR_WIDTH = 32,
    parameter HQM_SFI_RX_NDCRD = 4,
    parameter HQM_SFI_RX_NHCRD = 4,
    parameter HQM_SFI_RX_NUM_SHARED_POOLS = 0,
    parameter HQM_SFI_RX_PCIE_MERGED_SELECT = 0,
    parameter HQM_SFI_RX_PCIE_SHARED_SELECT = 0,
    parameter HQM_SFI_RX_RBN = 3,
    parameter HQM_SFI_RX_SHARED_CREDIT_EN = 0,
    parameter HQM_SFI_RX_SH_DATA_CRD_BLK_SZ = 1,
    parameter HQM_SFI_RX_SH_HDR_CRD_BLK_SZ = 1,
    parameter HQM_SFI_RX_TBN = 1,
    parameter HQM_SFI_RX_TX_CRD_REG = 1,
    parameter HQM_SFI_RX_VIRAL_EN = 0,
    parameter HQM_SFI_RX_VR = 0,
    parameter HQM_SFI_RX_VT = 0,
    parameter HQM_SFI_TX_BCM_EN = 1,
    parameter HQM_SFI_TX_BLOCK_EARLY_VLD_EN = 1,
    parameter HQM_SFI_TX_D = 32,
    parameter HQM_SFI_TX_DATA_AUX_PARITY_EN = 1,
    parameter HQM_SFI_TX_DATA_CRD_GRAN = 4,
    parameter HQM_SFI_TX_DATA_INTERLEAVE = 0,
    parameter HQM_SFI_TX_DATA_LAYER_EN = 1,
    parameter HQM_SFI_TX_DATA_MAX_FC_VC = 1,
    parameter HQM_SFI_TX_DATA_PARITY_EN = 1,
    parameter HQM_SFI_TX_DATA_PASS_HDR = 0,
    parameter HQM_SFI_TX_DS = 1,
    parameter HQM_SFI_TX_ECRC_SUPPORT = 0,
    parameter HQM_SFI_TX_FATAL_EN = 0,
    parameter HQM_SFI_TX_FLIT_MODE_PREFIX_EN = 0,
    parameter HQM_SFI_TX_H = 32,
    parameter HQM_SFI_TX_HDR_DATA_SEP = 0,
    parameter HQM_SFI_TX_HDR_MAX_FC_VC = 1,
    parameter HQM_SFI_TX_HGRAN = 4,
    parameter HQM_SFI_TX_HPARITY = 1,
    parameter HQM_SFI_TX_IDE_SUPPORT = 0,
    parameter HQM_SFI_TX_M = 1,
    parameter HQM_SFI_TX_MAX_CRD_CNT_WIDTH = 12,
    parameter HQM_SFI_TX_MAX_HDR_WIDTH = 32,
    parameter HQM_SFI_TX_NDCRD = 4,
    parameter HQM_SFI_TX_NHCRD = 4,
    parameter HQM_SFI_TX_NUM_SHARED_POOLS = 0,
    parameter HQM_SFI_TX_PCIE_MERGED_SELECT = 0,
    parameter HQM_SFI_TX_PCIE_SHARED_SELECT = 0,
    parameter HQM_SFI_TX_RBN = 1,
    parameter HQM_SFI_TX_SHARED_CREDIT_EN = 0,
    parameter HQM_SFI_TX_SH_DATA_CRD_BLK_SZ = 1,
    parameter HQM_SFI_TX_SH_HDR_CRD_BLK_SZ = 1,
    parameter HQM_SFI_TX_TBN = 3,
    parameter HQM_SFI_TX_TX_CRD_REG = 1,
    parameter HQM_SFI_TX_VIRAL_EN = 0,
    parameter HQM_SFI_TX_VR = 0,
    parameter HQM_SFI_TX_VT = 0,
    parameter HQM_TRIGFABWIDTH = 4,
    parameter HQM_TRIGGER_WIDTH = 3  ) (
    input           par_logic_pgcb_fet_en_ack_b,
    output          hqm_clk_enable,
    output          hqm_clk_rptr_rst_b,
    output          hqm_clk_trunk,
    output          hqm_clk_ungate,
    output          hqm_gated_rst_b,
    output          hqm_proc_reset_done_sync_hqm,
    output          prim_clk_enable,
    output          prim_clk_ungate,
    // Ports for Interface dvp_apb4
    input   [31:0]  dvp_paddr,
    input           dvp_penable,
    input   [2:0]   dvp_pprot,
    input           dvp_psel,
    input   [3:0]   dvp_pstrb,
    input   [31:0]  dvp_pwdata,
    input           dvp_pwrite,
    output  [31:0]  dvp_prdata,
    output          dvp_pready,
    output          dvp_pslverr,
    // Ports for Interface dvp_ctf
    input   [(HQM_TRIGFABWIDTH-1):0] ftrig_fabric_in,
    input   [(HQM_TRIGFABWIDTH-1):0] ftrig_fabric_out_ack,
    output  [(HQM_TRIGFABWIDTH-1):0] atrig_fabric_in_ack,
    output  [(HQM_TRIGFABWIDTH-1):0] atrig_fabric_out,
    // Ports for Interface dvp_dsp_inside
    input   [7:0]   fdfx_debug_cap,
    input           fdfx_debug_cap_valid,
    input           fdfx_earlyboot_debug_exit,
    input           fdfx_policy_update,
    input   [7:0]   fdfx_security_policy,
    // Ports for Interface dvp_dtf
    input           fdtf_upstream_active,
    input           fdtf_upstream_credit,
    input           fdtf_upstream_sync,
    output  [(HQM_DTF_DATA_WIDTH-1):0] adtf_dnstream_data,
    output  [(HQM_DTF_HEADER_WIDTH-1):0] adtf_dnstream_header,
    output          adtf_dnstream_valid,
    // Ports for Interface dvp_dtf_clock
    input           fdtf_clk,
    input           fdtf_cry_clk,
    // Ports for Interface dvp_dtf_misc
    input   [1:0]   fdtf_fast_cnt_width,
    input   [7:0]   fdtf_packetizer_cid,
    input   [7:0]   fdtf_packetizer_mid,
    input           fdtf_survive_mode,
    // Ports for Interface dvp_dtf_reset
    input           fdtf_rst_b,
    // Ports for Interface iosf_sideband
    input           gpsb_mnpcup,
    input           gpsb_mpccup,
    input   [2:0]   gpsb_side_ism_fabric,
    input           gpsb_teom,
    input           gpsb_tnpput,
    input           gpsb_tparity,
    input   [(HQM_SBE_DATAWIDTH-1):0] gpsb_tpayload,
    input           gpsb_tpcput,
    output          gpsb_meom,
    output          gpsb_mnpput,
    output          gpsb_mparity,
    output  [(HQM_SBE_DATAWIDTH-1):0] gpsb_mpayload,
    output          gpsb_mpcput,
    output  [2:0]   gpsb_side_ism_agent,
    output          gpsb_tnpcup,
    output          gpsb_tpccup,
    // Ports for Interface iosf_sideband_clock
    input           side_clk,
    // Ports for Interface iosf_sideband_idstraps
    input   [15:0]  strap_hqm_do_serr_dstid,
    input   [15:0]  strap_hqm_err_sb_dstid,
    input   [15:0]  strap_hqm_gpsb_srcid,
    // Ports for Interface iosf_sideband_pok
    output          side_pok,
    // Ports for Interface iosf_sideband_power
    input           side_clkack,
    output          side_clkreq,
    // Ports for Interface iosf_sideband_reset
    input           side_rst_b,
    // Ports for Interface iosf_sideband_wake
    input           side_pwrgate_pmc_wake,
    // Ports for Interface prim_clock_req_ack
    input           prim_clkack,
    output          prim_clkreq,
    // Ports for Interface prim_reset
    input           pma_safemode,
    input           powergood_rst_b,
    input           prim_pwrgate_pmc_wake,
    input           prim_rst_b,
    // Ports for Interface rtdr_iosfsb_ism
    input           rtdr_iosfsb_ism_capturedr,
    input           rtdr_iosfsb_ism_irdec,
    input           rtdr_iosfsb_ism_shiftdr,
    input           rtdr_iosfsb_ism_tdi,
    input           rtdr_iosfsb_ism_updatedr,
    output          rtdr_iosfsb_ism_tdo,
    // Ports for Interface rtdr_iosfsb_ism_clock
    input           rtdr_iosfsb_ism_tck,
    // Ports for Interface rtdr_iosfsb_ism_reset
    input           rtdr_iosfsb_ism_trst_b,
    // Ports for Interface rtdr_tapconfig
    input           rtdr_tapconfig_capturedr,
    input           rtdr_tapconfig_irdec,
    input           rtdr_tapconfig_shiftdr,
    input           rtdr_tapconfig_tdi,
    input           rtdr_tapconfig_updatedr,
    output          rtdr_tapconfig_tdo,
    // Ports for Interface rtdr_tapconfig_clock
    input           rtdr_tapconfig_tck,
    // Ports for Interface rtdr_tapconfig_reset
    input           rtdr_tapconfig_trst_b,
    // Ports for Interface rtdr_taptrigger
    input           rtdr_taptrigger_capturedr,
    input           rtdr_taptrigger_irdec,
    input           rtdr_taptrigger_shiftdr,
    input           rtdr_taptrigger_tdi,
    input           rtdr_taptrigger_updatedr,
    output          rtdr_taptrigger_tdo,
    // Ports for Interface rtdr_taptrigger_clock
    input           rtdr_taptrigger_tck,
    // Ports for Interface rtdr_taptrigger_reset
    input           rtdr_taptrigger_trst_b,
    // Ports for Interface scan
    input           fscan_byprst_b,
    input           fscan_clkungate,
    input           fscan_clkungate_syn,
    input           fscan_latchclosed_b,
    input           fscan_latchopen,
    input           fscan_mode,
    input           fscan_rstbypen,
    input           fscan_shiften,
    // Ports for Interface scan_reset
    input           fdfx_powergood,
    // Ports for Interface sfi_rx_data
    input   [((HQM_SFI_RX_D*8)-1):0] sfi_rx_data,
    input           sfi_rx_data_aux_parity,
    input           sfi_rx_data_crd_rtn_block,
    input           sfi_rx_data_early_valid,
    input   [((HQM_SFI_RX_D/4)-1):0] sfi_rx_data_edb,
    input   [((HQM_SFI_RX_D/4)-1):0] sfi_rx_data_end,
    input   [((HQM_SFI_RX_DS*8)-1):0] sfi_rx_data_info_byte,
    input   [((HQM_SFI_RX_D/8)-1):0] sfi_rx_data_parity,
    input   [((HQM_SFI_RX_D/4)-1):0] sfi_rx_data_poison,
    input           sfi_rx_data_start,
    input           sfi_rx_data_valid,
    output          sfi_rx_data_block,
    output  [1:0]   sfi_rx_data_crd_rtn_fc_id,
    output          sfi_rx_data_crd_rtn_valid,
    output  [(HQM_SFI_RX_NDCRD-1):0] sfi_rx_data_crd_rtn_value,
    output  [4:0]   sfi_rx_data_crd_rtn_vc_id,
    // Ports for Interface sfi_rx_globals
    input           sfi_rx_txcon_req,
    output          sfi_rx_rx_empty,
    output          sfi_rx_rxcon_ack,
    output          sfi_rx_rxdiscon_nack,
    // Ports for Interface sfi_rx_header
    input           sfi_rx_hdr_crd_rtn_block,
    input           sfi_rx_hdr_early_valid,
    input   [((HQM_SFI_RX_M*16)-1):0] sfi_rx_hdr_info_bytes,
    input           sfi_rx_hdr_valid,
    input   [((HQM_SFI_RX_H*8)-1):0] sfi_rx_header,
    output          sfi_rx_hdr_block,
    output  [1:0]   sfi_rx_hdr_crd_rtn_fc_id,
    output          sfi_rx_hdr_crd_rtn_valid,
    output  [(HQM_SFI_RX_NHCRD-1):0] sfi_rx_hdr_crd_rtn_value,
    output  [4:0]   sfi_rx_hdr_crd_rtn_vc_id,
    // Ports for Interface sfi_tx_data
    input           sfi_tx_data_block,
    input   [1:0]   sfi_tx_data_crd_rtn_fc_id,
    input           sfi_tx_data_crd_rtn_valid,
    input   [(HQM_SFI_TX_NDCRD-1):0] sfi_tx_data_crd_rtn_value,
    input   [4:0]   sfi_tx_data_crd_rtn_vc_id,
    output  [((HQM_SFI_TX_D*8)-1):0] sfi_tx_data,
    output          sfi_tx_data_aux_parity,
    output          sfi_tx_data_crd_rtn_block,
    output          sfi_tx_data_early_valid,
    output  [((HQM_SFI_TX_D/4)-1):0] sfi_tx_data_edb,
    output  [((HQM_SFI_TX_D/4)-1):0] sfi_tx_data_end,
    output  [((HQM_SFI_TX_DS*8)-1):0] sfi_tx_data_info_byte,
    output  [((HQM_SFI_TX_D/8)-1):0] sfi_tx_data_parity,
    output  [((HQM_SFI_TX_D/4)-1):0] sfi_tx_data_poison,
    output          sfi_tx_data_start,
    output          sfi_tx_data_valid,
    // Ports for Interface sfi_tx_globals
    input           sfi_tx_rx_empty,
    input           sfi_tx_rxcon_ack,
    input           sfi_tx_rxdiscon_nack,
    output          sfi_tx_txcon_req,
    // Ports for Interface sfi_tx_header
    input           sfi_tx_hdr_block,
    input   [1:0]   sfi_tx_hdr_crd_rtn_fc_id,
    input           sfi_tx_hdr_crd_rtn_valid,
    input   [(HQM_SFI_TX_NHCRD-1):0] sfi_tx_hdr_crd_rtn_value,
    input   [4:0]   sfi_tx_hdr_crd_rtn_vc_id,
    output          sfi_tx_hdr_crd_rtn_block,
    output          sfi_tx_hdr_early_valid,
    output  [((HQM_SFI_TX_M*16)-1):0] sfi_tx_hdr_info_bytes,
    output          sfi_tx_hdr_valid,
    output  [((HQM_SFI_TX_H*8)-1):0] sfi_tx_header,
    // Ports for Interface viewpins_dig
    output          dig_view_out_0,
    output          dig_view_out_1,
    // Ports for Manually exported pins
    input           ap_alarm_down_v,
    input           ap_alarm_up_ready,
    input           ap_aqed_ready,
    input           ap_aqed_v,
    input           ap_cfg_req_down_read,
    input           ap_cfg_req_down_write,
    input           ap_cfg_rsp_down_ack,
    input           ap_reset_done,
    input           ap_unit_idle,
    input           ap_unit_pipeidle,
    input           aqed_alarm_down_v,
    input           aqed_ap_enq_ready,
    input           aqed_ap_enq_v,
    input   [92:0]  aqed_cfg_req_down,
    input           aqed_cfg_req_down_read,
    input           aqed_cfg_req_down_write,
    input   [38:0]  aqed_cfg_rsp_down,
    input           aqed_cfg_rsp_down_ack,
    input           aqed_chp_sch_ready,
    input           aqed_chp_sch_v,
    input           aqed_lsp_sch_ready,
    input           aqed_lsp_sch_v,
    input           aqed_reset_done,
    input           aqed_unit_idle,
    input           aqed_unit_pipeidle,
    input           chp_alarm_up_ready,
    input           chp_cfg_req_down_read,
    input           chp_cfg_req_down_write,
    input           chp_cfg_rsp_down_ack,
    input           chp_lsp_cmp_ready,
    input           chp_lsp_cmp_v,
    input           chp_lsp_token_ready,
    input           chp_lsp_token_v,
    input           chp_reset_done,
    input           chp_rop_hcw_ready,
    input           chp_rop_hcw_v,
    input           chp_unit_idle,
    input           chp_unit_pipeidle,
    input           cwdi_interrupt_w_req_ready,
    input           cwdi_interrupt_w_req_valid,
    input           dp_lsp_enq_dir_ready,
    input           dp_lsp_enq_dir_v,
    input           dp_lsp_enq_rorply_ready,
    input           dp_lsp_enq_rorply_v,
    input           dp_reset_done,
    input           dp_unit_idle,
    input           dp_unit_pipeidle,
    input   [15:0]  early_fuses,
    input           fdfx_sbparity_def,
    input           fdtf_force_ts,
    input           fdtf_serial_download_tsc,
    input           fdtf_timestamp_valid,
    input   [55:0]  fdtf_timestamp_value,
    input   [15:0]  fdtf_tsc_adjustment_strap,
    input           hcw_enq_in_ready,
    input           hcw_enq_w_req_ready,
    input           hcw_enq_w_req_valid,
    input           hcw_sched_w_req_ready,
    input           hcw_sched_w_req_valid,
    input           hqm_alarm_ready,
    input           hqm_alarm_v,
    input           hqm_proc_clk_en_chp,
    input           hqm_proc_clk_en_dir,
    input           hqm_proc_clk_en_lsp,
    input           hqm_proc_clk_en_nalb,
    input           hqm_proc_clk_en_qed,
    input           hqm_proc_clk_en_sys,
    input   [29:0]  hqm_system_visa_str,
    input           i_hqm_AW_fet_en_sequencer_par_mem_pgcb_fet_en_ack_b,
    input           i_hqm_master_fscan_isol_ctrl,
    input           i_hqm_master_fscan_isol_lat_ctrl,
    input           i_hqm_master_fscan_ret_ctrl,
    input   [65:0]  i_hqm_sif_rf_ibcpl_data_fifo_rdata,
    input   [19:0]  i_hqm_sif_rf_ibcpl_hdr_fifo_rdata,
    input   [128:0] i_hqm_sif_rf_mstr_ll_data0_rdata,
    input   [128:0] i_hqm_sif_rf_mstr_ll_data1_rdata,
    input   [128:0] i_hqm_sif_rf_mstr_ll_data2_rdata,
    input   [128:0] i_hqm_sif_rf_mstr_ll_data3_rdata,
    input   [152:0] i_hqm_sif_rf_mstr_ll_hdr_rdata,
    input   [34:0]  i_hqm_sif_rf_mstr_ll_hpa_rdata,
    input   [32:0]  i_hqm_sif_rf_ri_tlq_fifo_npdata_rdata,
    input   [157:0] i_hqm_sif_rf_ri_tlq_fifo_nphdr_rdata,
    input   [263:0] i_hqm_sif_rf_ri_tlq_fifo_pdata_rdata,
    input   [152:0] i_hqm_sif_rf_ri_tlq_fifo_phdr_rdata,
    input   [9:0]   i_hqm_sif_rf_scrbd_mem_rdata,
    input   [38:0]  i_hqm_sif_rf_tlb_data0_4k_rdata,
    input   [38:0]  i_hqm_sif_rf_tlb_data1_4k_rdata,
    input   [38:0]  i_hqm_sif_rf_tlb_data2_4k_rdata,
    input   [38:0]  i_hqm_sif_rf_tlb_data3_4k_rdata,
    input   [38:0]  i_hqm_sif_rf_tlb_data4_4k_rdata,
    input   [38:0]  i_hqm_sif_rf_tlb_data5_4k_rdata,
    input   [38:0]  i_hqm_sif_rf_tlb_data6_4k_rdata,
    input   [38:0]  i_hqm_sif_rf_tlb_data7_4k_rdata,
    input   [84:0]  i_hqm_sif_rf_tlb_tag0_4k_rdata,
    input   [84:0]  i_hqm_sif_rf_tlb_tag1_4k_rdata,
    input   [84:0]  i_hqm_sif_rf_tlb_tag2_4k_rdata,
    input   [84:0]  i_hqm_sif_rf_tlb_tag3_4k_rdata,
    input   [84:0]  i_hqm_sif_rf_tlb_tag4_4k_rdata,
    input   [84:0]  i_hqm_sif_rf_tlb_tag5_4k_rdata,
    input   [84:0]  i_hqm_sif_rf_tlb_tag6_4k_rdata,
    input   [84:0]  i_hqm_sif_rf_tlb_tag7_4k_rdata,
    input   [1:0]   i_hqm_visa_hqm_core_visa_str_175_174,
    input   [1:0]   i_hqm_visa_hqm_core_visa_str_178_177,
    input   [1:0]   i_hqm_visa_hqm_core_visa_str_182_181,
    input   [1:0]   i_hqm_visa_hqm_core_visa_str_185_184,
    input   [1:0]   i_hqm_visa_hqm_core_visa_str_189_188,
    input   [1:0]   i_hqm_visa_hqm_core_visa_str_192_191,
    input   [1:0]   i_hqm_visa_hqm_core_visa_str_196_195,
    input   [1:0]   i_hqm_visa_hqm_core_visa_str_199_198,
    input   [1:0]   i_hqm_visa_hqm_core_visa_str_210_209,
    input   [1:0]   i_hqm_visa_hqm_core_visa_str_213_212,
    input   [1:0]   i_hqm_visa_hqm_core_visa_str_224_223,
    input   [1:0]   i_hqm_visa_hqm_core_visa_str_227_226,
    input   [1:0]   i_hqm_visa_hqm_core_visa_str_238_237,
    input   [1:0]   i_hqm_visa_hqm_core_visa_str_241_240,
    input           i_hqm_visa_hqm_core_visa_str_252,
    input           i_hqm_visa_hqm_core_visa_str_253,
    input           interrupt_w_req_ready,
    input           interrupt_w_req_valid,
    input           iosf_pgcb_clk,
    input           lsp_alarm_down_v,
    input           lsp_alarm_up_ready,
    input           lsp_cfg_req_down_read,
    input           lsp_cfg_req_down_write,
    input           lsp_cfg_rsp_down_ack,
    input           lsp_dp_sch_dir_ready,
    input           lsp_dp_sch_dir_v,
    input           lsp_dp_sch_rorply_ready,
    input           lsp_dp_sch_rorply_v,
    input           lsp_nalb_sch_atq_ready,
    input           lsp_nalb_sch_atq_v,
    input           lsp_nalb_sch_rorply_ready,
    input           lsp_nalb_sch_rorply_v,
    input           lsp_nalb_sch_unoord_ready,
    input           lsp_nalb_sch_unoord_v,
    input           lsp_reset_done,
    input           lsp_unit_idle,
    input           lsp_unit_pipeidle,
    input           nalb_lsp_enq_lb_ready,
    input           nalb_lsp_enq_lb_v,
    input           nalb_lsp_enq_rorply_ready,
    input           nalb_lsp_enq_rorply_v,
    input           nalb_reset_done,
    input           nalb_unit_idle,
    input           nalb_unit_pipeidle,
    input           pgcb_clk,
    input           pgcb_tck,
    input           pm_hqm_adr_assert,
    input           prim_clk,
    input           prochot,
    input           qed_alarm_down_v,
    input           qed_alarm_up_ready,
    input           qed_aqed_enq_ready,
    input           qed_aqed_enq_v,
    input           qed_cfg_req_down_read,
    input           qed_cfg_req_down_write,
    input           qed_cfg_rsp_down_ack,
    input           qed_chp_sch_ready,
    input           qed_chp_sch_v,
    input           qed_reset_done,
    input           qed_unit_idle,
    input           qed_unit_pipeidle,
    input           rop_alarm_down_v,
    input           rop_alarm_up_ready,
    input           rop_cfg_req_down_read,
    input           rop_cfg_req_down_write,
    input           rop_cfg_rsp_down_ack,
    input           rop_dp_enq_ready,
    input           rop_dp_enq_v,
    input           rop_dqed_enq_ready,
    input           rop_lsp_reordercmp_ready,
    input           rop_lsp_reordercmp_v,
    input           rop_nalb_enq_ready,
    input           rop_nalb_enq_v,
    input           rop_qed_dqed_enq_v,
    input           rop_qed_enq_ready,
    input           rop_qed_force_clockon,
    input           rop_reset_done,
    input           rop_unit_idle,
    input           rop_unit_pipeidle,
    input           sif_alarm_ready,
    input           strap_hqm_16b_portids,
    input   [7:0]   strap_hqm_cmpl_sai,
    input   [63:0]  strap_hqm_csr_cp,
    input   [63:0]  strap_hqm_csr_rac,
    input   [63:0]  strap_hqm_csr_wac,
    input   [15:0]  strap_hqm_device_id,
    input           strap_hqm_do_serr_rs,
    input   [7:0]   strap_hqm_do_serr_sai,
    input           strap_hqm_do_serr_sairs_valid,
    input   [2:0]   strap_hqm_do_serr_tag,
    input   [7:0]   strap_hqm_err_sb_sai,
    input   [7:0]   strap_hqm_force_pok_sai_0,
    input   [7:0]   strap_hqm_force_pok_sai_1,
    input   [7:0]   strap_hqm_resetprep_ack_sai,
    input   [7:0]   strap_hqm_resetprep_sai_0,
    input   [7:0]   strap_hqm_resetprep_sai_1,
    input   [7:0]   strap_hqm_tx_sai,
    input           strap_no_mgmt_acks,
    input           system_cfg_req_down_read,
    input           system_cfg_req_down_write,
    input           system_cfg_rsp_down_ack,
    input           system_idle,
    input           system_reset_done,
    input           visa_str_chp_lsp_cmp_data,
    input           wd_clkreq,
    input   [638:0] write_buffer_mstr,
    input           write_buffer_mstr_v,
    output  [160:0] hcw_enq_in_data,
    output          hcw_enq_in_v,
    output          hqm_flr_prep,
    output          hqm_gated_local_override,
    output          hqm_pm_adr_ack,
    output          i_hqm_AW_fet_en_sequencer_par_mem_pgcb_fet_en_b,
    output          i_hqm_master_pgcb_isol_en,
    output          i_hqm_master_pgcb_isol_en_b,
    output          i_hqm_pwrgood_rst_b_buf_o,
    output  [7:0]   i_hqm_sif_rf_ibcpl_data_fifo_raddr,
    output          i_hqm_sif_rf_ibcpl_data_fifo_rclk,
    output          i_hqm_sif_rf_ibcpl_data_fifo_rclk_rst_n,
    output          i_hqm_sif_rf_ibcpl_data_fifo_re,
    output  [7:0]   i_hqm_sif_rf_ibcpl_data_fifo_waddr,
    output          i_hqm_sif_rf_ibcpl_data_fifo_wclk,
    output          i_hqm_sif_rf_ibcpl_data_fifo_wclk_rst_n,
    output  [65:0]  i_hqm_sif_rf_ibcpl_data_fifo_wdata,
    output          i_hqm_sif_rf_ibcpl_data_fifo_we,
    output  [7:0]   i_hqm_sif_rf_ibcpl_hdr_fifo_raddr,
    output          i_hqm_sif_rf_ibcpl_hdr_fifo_rclk,
    output          i_hqm_sif_rf_ibcpl_hdr_fifo_rclk_rst_n,
    output          i_hqm_sif_rf_ibcpl_hdr_fifo_re,
    output  [7:0]   i_hqm_sif_rf_ibcpl_hdr_fifo_waddr,
    output          i_hqm_sif_rf_ibcpl_hdr_fifo_wclk,
    output          i_hqm_sif_rf_ibcpl_hdr_fifo_wclk_rst_n,
    output  [19:0]  i_hqm_sif_rf_ibcpl_hdr_fifo_wdata,
    output          i_hqm_sif_rf_ibcpl_hdr_fifo_we,
    output  [7:0]   i_hqm_sif_rf_mstr_ll_data0_raddr,
    output          i_hqm_sif_rf_mstr_ll_data0_rclk,
    output          i_hqm_sif_rf_mstr_ll_data0_rclk_rst_n,
    output          i_hqm_sif_rf_mstr_ll_data0_re,
    output  [7:0]   i_hqm_sif_rf_mstr_ll_data0_waddr,
    output          i_hqm_sif_rf_mstr_ll_data0_wclk,
    output          i_hqm_sif_rf_mstr_ll_data0_wclk_rst_n,
    output  [128:0] i_hqm_sif_rf_mstr_ll_data0_wdata,
    output          i_hqm_sif_rf_mstr_ll_data0_we,
    output  [7:0]   i_hqm_sif_rf_mstr_ll_data1_raddr,
    output          i_hqm_sif_rf_mstr_ll_data1_rclk,
    output          i_hqm_sif_rf_mstr_ll_data1_rclk_rst_n,
    output          i_hqm_sif_rf_mstr_ll_data1_re,
    output  [7:0]   i_hqm_sif_rf_mstr_ll_data1_waddr,
    output          i_hqm_sif_rf_mstr_ll_data1_wclk,
    output          i_hqm_sif_rf_mstr_ll_data1_wclk_rst_n,
    output  [128:0] i_hqm_sif_rf_mstr_ll_data1_wdata,
    output          i_hqm_sif_rf_mstr_ll_data1_we,
    output  [7:0]   i_hqm_sif_rf_mstr_ll_data2_raddr,
    output          i_hqm_sif_rf_mstr_ll_data2_rclk,
    output          i_hqm_sif_rf_mstr_ll_data2_rclk_rst_n,
    output          i_hqm_sif_rf_mstr_ll_data2_re,
    output  [7:0]   i_hqm_sif_rf_mstr_ll_data2_waddr,
    output          i_hqm_sif_rf_mstr_ll_data2_wclk,
    output          i_hqm_sif_rf_mstr_ll_data2_wclk_rst_n,
    output  [128:0] i_hqm_sif_rf_mstr_ll_data2_wdata,
    output          i_hqm_sif_rf_mstr_ll_data2_we,
    output  [7:0]   i_hqm_sif_rf_mstr_ll_data3_raddr,
    output          i_hqm_sif_rf_mstr_ll_data3_rclk,
    output          i_hqm_sif_rf_mstr_ll_data3_rclk_rst_n,
    output          i_hqm_sif_rf_mstr_ll_data3_re,
    output  [7:0]   i_hqm_sif_rf_mstr_ll_data3_waddr,
    output          i_hqm_sif_rf_mstr_ll_data3_wclk,
    output          i_hqm_sif_rf_mstr_ll_data3_wclk_rst_n,
    output  [128:0] i_hqm_sif_rf_mstr_ll_data3_wdata,
    output          i_hqm_sif_rf_mstr_ll_data3_we,
    output  [7:0]   i_hqm_sif_rf_mstr_ll_hdr_raddr,
    output          i_hqm_sif_rf_mstr_ll_hdr_rclk,
    output          i_hqm_sif_rf_mstr_ll_hdr_rclk_rst_n,
    output          i_hqm_sif_rf_mstr_ll_hdr_re,
    output  [7:0]   i_hqm_sif_rf_mstr_ll_hdr_waddr,
    output          i_hqm_sif_rf_mstr_ll_hdr_wclk,
    output          i_hqm_sif_rf_mstr_ll_hdr_wclk_rst_n,
    output  [152:0] i_hqm_sif_rf_mstr_ll_hdr_wdata,
    output          i_hqm_sif_rf_mstr_ll_hdr_we,
    output  [6:0]   i_hqm_sif_rf_mstr_ll_hpa_raddr,
    output          i_hqm_sif_rf_mstr_ll_hpa_rclk,
    output          i_hqm_sif_rf_mstr_ll_hpa_rclk_rst_n,
    output          i_hqm_sif_rf_mstr_ll_hpa_re,
    output  [6:0]   i_hqm_sif_rf_mstr_ll_hpa_waddr,
    output          i_hqm_sif_rf_mstr_ll_hpa_wclk,
    output          i_hqm_sif_rf_mstr_ll_hpa_wclk_rst_n,
    output  [34:0]  i_hqm_sif_rf_mstr_ll_hpa_wdata,
    output          i_hqm_sif_rf_mstr_ll_hpa_we,
    output  [2:0]   i_hqm_sif_rf_ri_tlq_fifo_npdata_raddr,
    output          i_hqm_sif_rf_ri_tlq_fifo_npdata_rclk,
    output          i_hqm_sif_rf_ri_tlq_fifo_npdata_rclk_rst_n,
    output          i_hqm_sif_rf_ri_tlq_fifo_npdata_re,
    output  [2:0]   i_hqm_sif_rf_ri_tlq_fifo_npdata_waddr,
    output          i_hqm_sif_rf_ri_tlq_fifo_npdata_wclk,
    output          i_hqm_sif_rf_ri_tlq_fifo_npdata_wclk_rst_n,
    output  [32:0]  i_hqm_sif_rf_ri_tlq_fifo_npdata_wdata,
    output          i_hqm_sif_rf_ri_tlq_fifo_npdata_we,
    output  [2:0]   i_hqm_sif_rf_ri_tlq_fifo_nphdr_raddr,
    output          i_hqm_sif_rf_ri_tlq_fifo_nphdr_rclk,
    output          i_hqm_sif_rf_ri_tlq_fifo_nphdr_rclk_rst_n,
    output          i_hqm_sif_rf_ri_tlq_fifo_nphdr_re,
    output  [2:0]   i_hqm_sif_rf_ri_tlq_fifo_nphdr_waddr,
    output          i_hqm_sif_rf_ri_tlq_fifo_nphdr_wclk,
    output          i_hqm_sif_rf_ri_tlq_fifo_nphdr_wclk_rst_n,
    output  [157:0] i_hqm_sif_rf_ri_tlq_fifo_nphdr_wdata,
    output          i_hqm_sif_rf_ri_tlq_fifo_nphdr_we,
    output  [4:0]   i_hqm_sif_rf_ri_tlq_fifo_pdata_raddr,
    output          i_hqm_sif_rf_ri_tlq_fifo_pdata_rclk,
    output          i_hqm_sif_rf_ri_tlq_fifo_pdata_rclk_rst_n,
    output          i_hqm_sif_rf_ri_tlq_fifo_pdata_re,
    output  [4:0]   i_hqm_sif_rf_ri_tlq_fifo_pdata_waddr,
    output          i_hqm_sif_rf_ri_tlq_fifo_pdata_wclk,
    output          i_hqm_sif_rf_ri_tlq_fifo_pdata_wclk_rst_n,
    output  [263:0] i_hqm_sif_rf_ri_tlq_fifo_pdata_wdata,
    output          i_hqm_sif_rf_ri_tlq_fifo_pdata_we,
    output  [3:0]   i_hqm_sif_rf_ri_tlq_fifo_phdr_raddr,
    output          i_hqm_sif_rf_ri_tlq_fifo_phdr_rclk,
    output          i_hqm_sif_rf_ri_tlq_fifo_phdr_rclk_rst_n,
    output          i_hqm_sif_rf_ri_tlq_fifo_phdr_re,
    output  [3:0]   i_hqm_sif_rf_ri_tlq_fifo_phdr_waddr,
    output          i_hqm_sif_rf_ri_tlq_fifo_phdr_wclk,
    output          i_hqm_sif_rf_ri_tlq_fifo_phdr_wclk_rst_n,
    output  [152:0] i_hqm_sif_rf_ri_tlq_fifo_phdr_wdata,
    output          i_hqm_sif_rf_ri_tlq_fifo_phdr_we,
    output  [7:0]   i_hqm_sif_rf_scrbd_mem_raddr,
    output          i_hqm_sif_rf_scrbd_mem_rclk,
    output          i_hqm_sif_rf_scrbd_mem_rclk_rst_n,
    output          i_hqm_sif_rf_scrbd_mem_re,
    output  [7:0]   i_hqm_sif_rf_scrbd_mem_waddr,
    output          i_hqm_sif_rf_scrbd_mem_wclk,
    output          i_hqm_sif_rf_scrbd_mem_wclk_rst_n,
    output  [9:0]   i_hqm_sif_rf_scrbd_mem_wdata,
    output          i_hqm_sif_rf_scrbd_mem_we,
    output  [3:0]   i_hqm_sif_rf_tlb_data0_4k_raddr,
    output          i_hqm_sif_rf_tlb_data0_4k_rclk,
    output          i_hqm_sif_rf_tlb_data0_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_data0_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_data0_4k_waddr,
    output          i_hqm_sif_rf_tlb_data0_4k_wclk,
    output          i_hqm_sif_rf_tlb_data0_4k_wclk_rst_n,
    output  [38:0]  i_hqm_sif_rf_tlb_data0_4k_wdata,
    output          i_hqm_sif_rf_tlb_data0_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_data1_4k_raddr,
    output          i_hqm_sif_rf_tlb_data1_4k_rclk,
    output          i_hqm_sif_rf_tlb_data1_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_data1_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_data1_4k_waddr,
    output          i_hqm_sif_rf_tlb_data1_4k_wclk,
    output          i_hqm_sif_rf_tlb_data1_4k_wclk_rst_n,
    output  [38:0]  i_hqm_sif_rf_tlb_data1_4k_wdata,
    output          i_hqm_sif_rf_tlb_data1_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_data2_4k_raddr,
    output          i_hqm_sif_rf_tlb_data2_4k_rclk,
    output          i_hqm_sif_rf_tlb_data2_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_data2_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_data2_4k_waddr,
    output          i_hqm_sif_rf_tlb_data2_4k_wclk,
    output          i_hqm_sif_rf_tlb_data2_4k_wclk_rst_n,
    output  [38:0]  i_hqm_sif_rf_tlb_data2_4k_wdata,
    output          i_hqm_sif_rf_tlb_data2_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_data3_4k_raddr,
    output          i_hqm_sif_rf_tlb_data3_4k_rclk,
    output          i_hqm_sif_rf_tlb_data3_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_data3_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_data3_4k_waddr,
    output          i_hqm_sif_rf_tlb_data3_4k_wclk,
    output          i_hqm_sif_rf_tlb_data3_4k_wclk_rst_n,
    output  [38:0]  i_hqm_sif_rf_tlb_data3_4k_wdata,
    output          i_hqm_sif_rf_tlb_data3_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_data4_4k_raddr,
    output          i_hqm_sif_rf_tlb_data4_4k_rclk,
    output          i_hqm_sif_rf_tlb_data4_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_data4_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_data4_4k_waddr,
    output          i_hqm_sif_rf_tlb_data4_4k_wclk,
    output          i_hqm_sif_rf_tlb_data4_4k_wclk_rst_n,
    output  [38:0]  i_hqm_sif_rf_tlb_data4_4k_wdata,
    output          i_hqm_sif_rf_tlb_data4_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_data5_4k_raddr,
    output          i_hqm_sif_rf_tlb_data5_4k_rclk,
    output          i_hqm_sif_rf_tlb_data5_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_data5_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_data5_4k_waddr,
    output          i_hqm_sif_rf_tlb_data5_4k_wclk,
    output          i_hqm_sif_rf_tlb_data5_4k_wclk_rst_n,
    output  [38:0]  i_hqm_sif_rf_tlb_data5_4k_wdata,
    output          i_hqm_sif_rf_tlb_data5_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_data6_4k_raddr,
    output          i_hqm_sif_rf_tlb_data6_4k_rclk,
    output          i_hqm_sif_rf_tlb_data6_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_data6_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_data6_4k_waddr,
    output          i_hqm_sif_rf_tlb_data6_4k_wclk,
    output          i_hqm_sif_rf_tlb_data6_4k_wclk_rst_n,
    output  [38:0]  i_hqm_sif_rf_tlb_data6_4k_wdata,
    output          i_hqm_sif_rf_tlb_data6_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_data7_4k_raddr,
    output          i_hqm_sif_rf_tlb_data7_4k_rclk,
    output          i_hqm_sif_rf_tlb_data7_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_data7_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_data7_4k_waddr,
    output          i_hqm_sif_rf_tlb_data7_4k_wclk,
    output          i_hqm_sif_rf_tlb_data7_4k_wclk_rst_n,
    output  [38:0]  i_hqm_sif_rf_tlb_data7_4k_wdata,
    output          i_hqm_sif_rf_tlb_data7_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_tag0_4k_raddr,
    output          i_hqm_sif_rf_tlb_tag0_4k_rclk,
    output          i_hqm_sif_rf_tlb_tag0_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_tag0_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_tag0_4k_waddr,
    output          i_hqm_sif_rf_tlb_tag0_4k_wclk,
    output          i_hqm_sif_rf_tlb_tag0_4k_wclk_rst_n,
    output  [84:0]  i_hqm_sif_rf_tlb_tag0_4k_wdata,
    output          i_hqm_sif_rf_tlb_tag0_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_tag1_4k_raddr,
    output          i_hqm_sif_rf_tlb_tag1_4k_rclk,
    output          i_hqm_sif_rf_tlb_tag1_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_tag1_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_tag1_4k_waddr,
    output          i_hqm_sif_rf_tlb_tag1_4k_wclk,
    output          i_hqm_sif_rf_tlb_tag1_4k_wclk_rst_n,
    output  [84:0]  i_hqm_sif_rf_tlb_tag1_4k_wdata,
    output          i_hqm_sif_rf_tlb_tag1_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_tag2_4k_raddr,
    output          i_hqm_sif_rf_tlb_tag2_4k_rclk,
    output          i_hqm_sif_rf_tlb_tag2_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_tag2_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_tag2_4k_waddr,
    output          i_hqm_sif_rf_tlb_tag2_4k_wclk,
    output          i_hqm_sif_rf_tlb_tag2_4k_wclk_rst_n,
    output  [84:0]  i_hqm_sif_rf_tlb_tag2_4k_wdata,
    output          i_hqm_sif_rf_tlb_tag2_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_tag3_4k_raddr,
    output          i_hqm_sif_rf_tlb_tag3_4k_rclk,
    output          i_hqm_sif_rf_tlb_tag3_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_tag3_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_tag3_4k_waddr,
    output          i_hqm_sif_rf_tlb_tag3_4k_wclk,
    output          i_hqm_sif_rf_tlb_tag3_4k_wclk_rst_n,
    output  [84:0]  i_hqm_sif_rf_tlb_tag3_4k_wdata,
    output          i_hqm_sif_rf_tlb_tag3_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_tag4_4k_raddr,
    output          i_hqm_sif_rf_tlb_tag4_4k_rclk,
    output          i_hqm_sif_rf_tlb_tag4_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_tag4_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_tag4_4k_waddr,
    output          i_hqm_sif_rf_tlb_tag4_4k_wclk,
    output          i_hqm_sif_rf_tlb_tag4_4k_wclk_rst_n,
    output  [84:0]  i_hqm_sif_rf_tlb_tag4_4k_wdata,
    output          i_hqm_sif_rf_tlb_tag4_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_tag5_4k_raddr,
    output          i_hqm_sif_rf_tlb_tag5_4k_rclk,
    output          i_hqm_sif_rf_tlb_tag5_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_tag5_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_tag5_4k_waddr,
    output          i_hqm_sif_rf_tlb_tag5_4k_wclk,
    output          i_hqm_sif_rf_tlb_tag5_4k_wclk_rst_n,
    output  [84:0]  i_hqm_sif_rf_tlb_tag5_4k_wdata,
    output          i_hqm_sif_rf_tlb_tag5_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_tag6_4k_raddr,
    output          i_hqm_sif_rf_tlb_tag6_4k_rclk,
    output          i_hqm_sif_rf_tlb_tag6_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_tag6_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_tag6_4k_waddr,
    output          i_hqm_sif_rf_tlb_tag6_4k_wclk,
    output          i_hqm_sif_rf_tlb_tag6_4k_wclk_rst_n,
    output  [84:0]  i_hqm_sif_rf_tlb_tag6_4k_wdata,
    output          i_hqm_sif_rf_tlb_tag6_4k_we,
    output  [3:0]   i_hqm_sif_rf_tlb_tag7_4k_raddr,
    output          i_hqm_sif_rf_tlb_tag7_4k_rclk,
    output          i_hqm_sif_rf_tlb_tag7_4k_rclk_rst_n,
    output          i_hqm_sif_rf_tlb_tag7_4k_re,
    output  [3:0]   i_hqm_sif_rf_tlb_tag7_4k_waddr,
    output          i_hqm_sif_rf_tlb_tag7_4k_wclk,
    output          i_hqm_sif_rf_tlb_tag7_4k_wclk_rst_n,
    output  [84:0]  i_hqm_sif_rf_tlb_tag7_4k_wdata,
    output          i_hqm_sif_rf_tlb_tag7_4k_we,
    output          ip_ready,
    output          logic_pgcb_fet_en_b,
    output  [15:0]  master_chp_timestamp,
    output  [92:0]  mstr_cfg_req_down,
    output          mstr_cfg_req_down_read,
    output          mstr_cfg_req_down_write,
    output          pci_cfg_pmsixctl_fm,
    output          pci_cfg_pmsixctl_msie,
    output          pci_cfg_sciov_en,
    output          reset_prep_ack,
    output  [24:0]  sif_alarm_data,
    output          sif_alarm_v,
    output          write_buffer_mstr_ready
);

   wire         final_pgcb_fet_en_ack_b;
   wire         flr_triggered;
   wire         fuse_force_on;
   wire         fuse_proc_disable;
   wire         hqm_cdc_clk;
   wire         hqm_cdc_clk_enable_mstr;
   wire         hqm_cdc_clk_enable_rptr;
   wire [23:0]  hqm_cdc_visa;
   wire         hqm_clk_rptr_rst_sync_b;
   wire         hqm_clk_throttle;
   wire         hqm_clk_ungate_rptr;
   wire [0:0]   hqm_freerun_clk_enable_and_mstr;
   wire         hqm_freerun_clk_enable_rptr_mstr;
   wire         hqm_freerun_clk_mstr;
   wire         hqm_gated_rst_b_mstr;
   wire         hqm_gclock_enable;
   wire         hqm_inp_gated_clk;
   wire         hqm_inp_gated_clk_enable_rptr;
   wire [0:0]   hqm_master_hqm_cdc_enable;
   wire [23:0]  hqm_pgcb_visa;
   wire [31:0]  hqm_pmsm_visa;
   wire         hqm_proc_clkreq_b;
   wire         hqm_proc_reset_done;
   wire         hqm_pwrgood_rst_b_internal;
   wire         hqm_shields_up;
   wire [679:0] hqm_sif_visa;
   wire [9:0]   hqm_triggers_in;
   wire         i_hqm_master_hqm_cfg_master_clkreq_b;
   wire         i_hqm_master_hqm_clk_enable;
   wire         i_hqm_master_hqm_clk_rptr_rst_b;
   wire         i_hqm_master_hqm_clk_ungate;
   wire         i_hqm_master_hqm_proc_reset_done_sync_hqm;
   wire         i_hqm_master_pgcb_fet_en_b;
   wire         i_hqm_sif_prim_clk_enable;
   wire         i_hqm_sif_prim_clk_ungate;
   wire         i_system_buf_hqm_clk_trunk_o;
   wire [31:0]  master_ctl;
   wire         master_ctl_load;
   wire         nonflr_clk_enable_rptr;
   wire [31:0]  paddr;
   wire         penable;
   wire         pgcb_fet_en_ack_b;
   wire         pgcb_fet_en_b_out;
   wire         pgcb_force_rst_b;
   wire         pgcb_hqm_pwrgate_active;
   wire         pgcb_isol_en_b;
   wire         pm_allow_ing_drop;
   wire         pm_fsm_active;
   wire         pm_fsm_d0tod3_ok;
   wire         pm_fsm_d3tod0_ok;
   wire         pm_fsm_in_run;
   wire [1:0]   pm_state;
   wire [31:0]  prdata;
   wire         prdata_par;
   wire         pready;
   wire         prim_clk_enable_cdc;
   wire         prim_clk_enable_rptr;
   wire         prim_clk_enable_rptr_mstr;
   wire         prim_clk_enable_sys;
   wire         prim_clk_ungate_rptr;
   wire         prim_gated_clk;
   wire         prim_gated_clk_mstr;
   wire         prim_gated_rst_b;
   wire         prim_nonflr_clk;
   wire         psel;
   wire         pslverr;
   wire [19:0]  puser;
   wire [31:0]  pwdata;
   wire         pwrite;
   wire [31:0]  rtdr_func_po_iosfsb_ism;
   wire [31:0]  rtdr_func_po_tapconfig;
   wire [31:0]  rtdr_func_po_taptrigger;
   wire         side_rst_sync_prim_n;
   wire         visa_str_hqm_cdc_clk_enable;
   wire         visa_str_hqm_clk_enable;
   wire         visa_str_hqm_clk_throttle;
   wire         visa_str_hqm_flr_prep;
   wire         visa_str_hqm_gated_local_override;
   wire         visa_str_hqm_gclock_enable;
   wire         visa_str_hqm_proc_idle;
   wire         visa_str_hqm_proc_pipeidle;
   wire         visa_str_pm_ip_clk_halt_b_2_rpt_0_iosf;
   wire         visa_str_prim_clk_enable;

   hqm_AW_fet_en_sequencer i_hqm_AW_fet_en_sequencer
      (.pgcb_fet_en_b               (i_hqm_master_pgcb_fet_en_b),
       .par_logic_pgcb_fet_en_b     (logic_pgcb_fet_en_b),
       .par_mem_pgcb_fet_en_b       (i_hqm_AW_fet_en_sequencer_par_mem_pgcb_fet_en_b),
       .par_logic_pgcb_fet_en_ack_b,
       .par_mem_pgcb_fet_en_ack_b   (i_hqm_AW_fet_en_sequencer_par_mem_pgcb_fet_en_ack_b),
       .pgcb_fet_en_ack_b);

   hqm_AW_viewpin_mux
      #(.NUM_IN(7),
        .MUX_SEL_WIDTH(3),
        .NUM_OUT(2)) i_hqm_AW_viewpin_mux
      (.mux_in  ({pgcb_fet_en_b_out, 
                  final_pgcb_fet_en_ack_b, 
                  pgcb_hqm_pwrgate_active, 
                  pgcb_isol_en_b, 
                  pgcb_force_rst_b, 
                  pm_fsm_active, 
                  hqm_cdc_clk_enable_mstr}),
       .mux_sel (rtdr_func_po_tapconfig[10:5]),
       .mux_out ({dig_view_out_1, dig_view_out_0}));

   hqm_master
      #(.HQM_TRIGGER_WIDTH(HQM_TRIGGER_WIDTH)) i_hqm_master
      (.prim_gated_clk                         (prim_gated_clk_mstr),
       .prim_clk_enable                        (prim_clk_enable_rptr_mstr),
       .hqm_freerun_clk                        (hqm_freerun_clk_mstr),
       .hqm_fullrate_clk                       (i_system_buf_hqm_clk_trunk_o),
       .hqm_clk_ungate                         (i_hqm_master_hqm_clk_ungate),
       .hqm_clk_enable                         (i_hqm_master_hqm_clk_enable),
       .hqm_clk_throttle,
       .hqm_gclock_enable,
       .hqm_cdc_clk,
       .hqm_inp_gated_clk,
       .prim_freerun_clk                       (prim_clk),
       .aon_clk                                (fdtf_clk),
       .pgcb_clk,
       .wd_clkreq,
       .hqm_proc_clkreq_b,
       // Tie to constant value: one
       .pm_ip_clk_halt_b_2_rpt_0_iosf          (1'b1),
       .side_rst_b,
       .prim_gated_rst_b,
       .hqm_gated_rst_b                        (hqm_gated_rst_b_mstr),
       .hqm_clk_rptr_rst_b                     (i_hqm_master_hqm_clk_rptr_rst_b),
       .flr_triggered,
       .hqm_shields_up,
       .hqm_flr_prep,
       .hqm_pwrgood_rst_b                      (hqm_pwrgood_rst_b_internal),
       .hqm_gated_local_override,
       .prochot,
       .pm_state,
       .master_ctl_load,
       .master_ctl,
       .pm_fsm_d0tod3_ok,
       .pm_fsm_d3tod0_ok,
       .pm_fsm_in_run,
       .pm_allow_ing_drop,
       .pgcb_isol_en_b,
       .pgcb_isol_en                           (i_hqm_master_pgcb_isol_en),
       .pgcb_fet_en_b                          (i_hqm_master_pgcb_fet_en_b),
       .pgcb_fet_en_ack_b,
       .fuse_force_on,
       .fuse_proc_disable,
       .master_chp_timestamp,
       .puser,
       .psel,
       .pwrite,
       .penable,
       .paddr,
       .pwdata,
       .pready,
       .pslverr,
       .prdata,
       .prdata_par,
       .mstr_cfg_req_down_write,
       .mstr_cfg_req_down_read,
       .mstr_cfg_req_down,
       .mstr_cfg_rsp_up_ack                    (aqed_cfg_rsp_down_ack),
       .mstr_cfg_rsp_up                        (aqed_cfg_rsp_down),
       .mstr_cfg_req_up_write                  (aqed_cfg_req_down_write),
       .mstr_cfg_req_up_read                   (aqed_cfg_req_down_read),
       .mstr_cfg_req_up                        (aqed_cfg_req_down),
       .mstr_hqm_reset_done                    ({system_reset_done, 
                                                 aqed_reset_done, 
                                                 qed_reset_done, 
                                                 qed_reset_done, 
                                                 dp_reset_done, 
                                                 ap_reset_done, 
                                                 nalb_reset_done, 
                                                 lsp_reset_done, 
                                                 rop_reset_done, 
                                                 chp_reset_done}),
       .mstr_unit_idle                         ({system_idle, 
                                                 aqed_unit_idle, 
                                                 qed_unit_idle, 
                                                 qed_unit_idle, 
                                                 dp_unit_idle, 
                                                 ap_unit_idle, 
                                                 nalb_unit_idle, 
                                                 lsp_unit_idle, 
                                                 rop_unit_idle, 
                                                 chp_unit_idle}),
       // Tie to constant value: one
       .mstr_unit_pipeidle                     ({1'b1, 
                                                 aqed_unit_pipeidle, 
                                                 qed_unit_pipeidle, 
                                                 qed_unit_pipeidle, 
                                                 dp_unit_pipeidle, 
                                                 ap_unit_pipeidle, 
                                                 nalb_unit_pipeidle, 
                                                 lsp_unit_pipeidle, 
                                                 rop_unit_pipeidle, 
                                                 chp_unit_pipeidle}),
       .mstr_lcb_enable                        ({hqm_proc_clk_en_sys, 
                                                 hqm_proc_clk_en_lsp, 
                                                 hqm_proc_clk_en_qed, 
                                                 hqm_proc_clk_en_qed, 
                                                 hqm_proc_clk_en_nalb, 
                                                 hqm_proc_clk_en_lsp, 
                                                 hqm_proc_clk_en_dir, 
                                                 hqm_proc_clk_en_lsp, 
                                                 hqm_proc_clk_en_chp, 
                                                 hqm_proc_clk_en_chp}),
       .hqm_proc_reset_done_sync_hqm           (i_hqm_master_hqm_proc_reset_done_sync_hqm),
       .hqm_proc_reset_done,
       .visa_str_hqm_proc_idle,
       .visa_str_hqm_proc_pipeidle,
       .visa_str_prim_clk_enable,
       .visa_str_hqm_clk_enable,
       .visa_str_hqm_clk_throttle,
       .visa_str_hqm_gclock_enable,
       .visa_str_hqm_cdc_clk_enable,
       .visa_str_hqm_gated_local_override,
       .visa_str_hqm_flr_prep,
       .visa_str_pm_ip_clk_halt_b_2_rpt_0_iosf,
       .hqm_triggers_in,
       .hqm_triggers                           (),
       .pgcb_tck,
       .fdfx_powergood,
       .fdfx_pgcb_bypass                       (rtdr_func_po_tapconfig[1]),
       .fdfx_pgcb_ovr                          (rtdr_func_po_tapconfig[2]),
       .fscan_ret_ctrl                         (i_hqm_master_fscan_ret_ctrl),
       .fscan_isol_ctrl                        (i_hqm_master_fscan_isol_ctrl),
       .fscan_isol_lat_ctrl                    (i_hqm_master_fscan_isol_lat_ctrl),
       .fscan_clkungate,
       .fscan_rstbypen,
       .fscan_byprst_b,
       .fscan_mode,
       .fscan_fet_on                           (rtdr_func_po_tapconfig[3]),
       .fscan_trigger_mask_v                   (rtdr_func_po_taptrigger[30]),
       .fscan_trigger_mask                     (rtdr_func_po_taptrigger[29:0]),
       .fscan_fet_en_sel                       (rtdr_func_po_tapconfig[4]),
       .cdc_hqm_jta_force_clkreq               (rtdr_func_po_iosfsb_ism[2]),
       .cdc_hqm_jta_clkgate_ovrd               (rtdr_func_po_iosfsb_ism[1]),
       .hqm_cdc_clk_enable                     (hqm_cdc_clk_enable_mstr),
       .hw_reset_force_pwr_on                  (rtdr_func_po_tapconfig[11]),
       .pgcb_hqm_pwrgate_active,
       .final_pgcb_fet_en_ack_b,
       .pgcb_fet_en_b_out,
       .pgcb_force_rst_b,
       .pm_fsm_active,
       .hqm_cdc_visa,
       .hqm_pgcbunit_visa                      (hqm_pgcb_visa),
       .hqm_pmsm_visa,
       .hqm_cfg_master_clkreq_b                (i_hqm_master_hqm_cfg_master_clkreq_b));

   hqm_AW_clkgate i_hqm_master_clkfree
      (.clk             (i_system_buf_hqm_clk_trunk_o),
       .enable          (hqm_freerun_clk_enable_rptr_mstr),
       .cfg_clkungate   (hqm_clk_ungate_rptr),
       .fscan_clkungate,
       .gated_clk       (hqm_freerun_clk_mstr));

   hqm_AW_flop i_hqm_master_hqm_cdc_clk_enable_rptr
      (.clk    (i_system_buf_hqm_clk_trunk_o),
       .rst_n  (hqm_clk_rptr_rst_sync_b),
       .data   (hqm_cdc_clk_enable_mstr),
       .data_q (hqm_cdc_clk_enable_rptr));

   hqm_AW_clkgate i_hqm_master_hqm_cdc_clkgate
      (.clk             (i_system_buf_hqm_clk_trunk_o),
       .enable          (hqm_master_hqm_cdc_enable),
       .cfg_clkungate   (hqm_clk_ungate_rptr),
       .fscan_clkungate,
       .gated_clk       (hqm_cdc_clk));

   hqm_AW_clkand2_comb
      #(.WIDTH(1)) i_hqm_master_hqm_cdc_enable_and2
      (.clki0 (hqm_cdc_clk_enable_rptr),
       .clki1 (hqm_clk_rptr_rst_sync_b),
       .clko  (hqm_master_hqm_cdc_enable));

   hqm_AW_reset_sync_scan i_hqm_master_hqm_clk_rptr_rst_sync_n
      (.clk            (i_system_buf_hqm_clk_trunk_o),
       .rst_n          (i_hqm_master_hqm_clk_rptr_rst_b),
       .fscan_rstbypen,
       .fscan_byprst_b,
       .rst_n_sync     (hqm_clk_rptr_rst_sync_b));

   hqm_AW_flop i_hqm_master_hqm_clk_ungate_rptr
      (.clk    (i_system_buf_hqm_clk_trunk_o),
       .rst_n  (hqm_clk_rptr_rst_sync_b),
       .data   (i_hqm_master_hqm_clk_ungate),
       .data_q (hqm_clk_ungate_rptr));

   hqm_AW_clkand2_comb
      #(.WIDTH(1)) i_hqm_master_hqm_freerun_clk_enable_and2
      (.clki0 (hqm_clk_throttle),
       .clki1 (hqm_gclock_enable),
       .clko  (hqm_freerun_clk_enable_and_mstr));

   hqm_AW_flop i_hqm_master_hqm_freerun_clk_enable_rptr
      (.clk    (i_system_buf_hqm_clk_trunk_o),
       .rst_n  (hqm_clk_rptr_rst_sync_b),
       .data   (hqm_freerun_clk_enable_and_mstr),
       .data_q (hqm_freerun_clk_enable_rptr_mstr));

   hqm_AW_clkgate i_hqm_master_hqm_inp_clkgate
      (.clk             (i_system_buf_hqm_clk_trunk_o),
       .enable          (hqm_inp_gated_clk_enable_rptr),
       .cfg_clkungate   (hqm_clk_ungate_rptr),
       .fscan_clkungate,
       .gated_clk       (hqm_inp_gated_clk));

   hqm_AW_flop i_hqm_master_hqm_inp_gated_clk_enable_rptr
      (.clk    (i_system_buf_hqm_clk_trunk_o),
       .rst_n  (hqm_clk_rptr_rst_sync_b),
       .data   (i_hqm_master_hqm_clk_enable),
       .data_q (hqm_inp_gated_clk_enable_rptr));

   hqm_AW_flop i_hqm_master_prim_clk_enable_rptr
      (.clk    (prim_clk),
       .rst_n  (side_rst_sync_prim_n),
       .data   (i_hqm_sif_prim_clk_enable),
       .data_q (prim_clk_enable_rptr_mstr));

   hqm_AW_flop i_hqm_master_prim_clk_ungate_rptr
      (.clk    (prim_clk),
       .rst_n  (side_rst_sync_prim_n),
       .data   (i_hqm_sif_prim_clk_ungate),
       .data_q (prim_clk_ungate_rptr));

   hqm_AW_clkgate i_hqm_master_prim_clkgate
      (.clk             (prim_clk),
       .enable          (prim_clk_enable_rptr_mstr),
       .cfg_clkungate   (prim_clk_ungate_rptr),
       .fscan_clkungate,
       .gated_clk       (prim_gated_clk_mstr));

   hqm_AW_reset_sync_scan i_hqm_master_side_rst_sync_prim_n
      (.clk            (prim_clk),
       .rst_n          (side_rst_b),
       .fscan_rstbypen,
       .fscan_byprst_b,
       .rst_n_sync     (side_rst_sync_prim_n));

   hqm_AW_buf i_hqm_pwrgood_rst_b_buf
      (.a (hqm_pwrgood_rst_b_internal),
       .o (i_hqm_pwrgood_rst_b_buf_o));

   hqm_AW_rtdr_reg
      #(.DWIDTH(32)) i_hqm_rtdr_iosfsb_ism
      (.tck       (rtdr_iosfsb_ism_tck),
       .trstb     (rtdr_iosfsb_ism_trst_b),
       .tdi       (rtdr_iosfsb_ism_tdi),
       .irdec     (rtdr_iosfsb_ism_irdec),
       .shiftdr   (rtdr_iosfsb_ism_shiftdr),
       .updatedr  (rtdr_iosfsb_ism_updatedr),
       .capturedr (rtdr_iosfsb_ism_capturedr),
       // Collage will use this name for the whole bus
       .func_pi   (rtdr_func_po_iosfsb_ism),
       .tdo       (rtdr_iosfsb_ism_tdo),
       // Collage will use this name for the whole bus
       .func_po   (rtdr_func_po_iosfsb_ism));

   hqm_AW_rtdr_reg
      #(.DWIDTH(32)) i_hqm_rtdr_tapconfig
      (.tck       (rtdr_tapconfig_tck),
       .trstb     (rtdr_tapconfig_trst_b),
       .tdi       (rtdr_tapconfig_tdi),
       .irdec     (rtdr_tapconfig_irdec),
       .shiftdr   (rtdr_tapconfig_shiftdr),
       .updatedr  (rtdr_tapconfig_updatedr),
       .capturedr (rtdr_tapconfig_capturedr),
       // Collage will use this name for the whole bus
       .func_pi   (rtdr_func_po_tapconfig),
       .tdo       (rtdr_tapconfig_tdo),
       // Collage will use this name for the whole bus
       .func_po   (rtdr_func_po_tapconfig));

   hqm_AW_rtdr_reg
      #(.DWIDTH(32)) i_hqm_rtdr_taptrigger
      (.tck       (rtdr_taptrigger_tck),
       .trstb     (rtdr_taptrigger_trst_b),
       .tdi       (rtdr_taptrigger_tdi),
       .irdec     (rtdr_taptrigger_irdec),
       .shiftdr   (rtdr_taptrigger_shiftdr),
       .updatedr  (rtdr_taptrigger_updatedr),
       .capturedr (rtdr_taptrigger_capturedr),
       // Collage wll use this name for the whole bus
       .func_pi   (rtdr_func_po_taptrigger),
       .tdo       (rtdr_taptrigger_tdo),
       // Collage wll use this name for the whole bus
       .func_po   (rtdr_func_po_taptrigger));

   hqm_sif
      #(.HQM_SBE_NPQUEUEDEPTH(HQM_SBE_NPQUEUEDEPTH),
        .HQM_SBE_PCQUEUEDEPTH(HQM_SBE_PCQUEUEDEPTH),
        .HQM_SBE_DATAWIDTH(HQM_SBE_DATAWIDTH),
        .HQM_SBE_PARITY_REQUIRED(HQM_SBE_PARITY_REQUIRED),
        .HQM_SFI_RX_BCM_EN(HQM_SFI_RX_BCM_EN),
        .HQM_SFI_RX_BLOCK_EARLY_VLD_EN(HQM_SFI_RX_BLOCK_EARLY_VLD_EN),
        .HQM_SFI_RX_D(HQM_SFI_RX_D),
        .HQM_SFI_RX_DATA_AUX_PARITY_EN(HQM_SFI_RX_DATA_AUX_PARITY_EN),
        .HQM_SFI_RX_DATA_CRD_GRAN(HQM_SFI_RX_DATA_CRD_GRAN),
        .HQM_SFI_RX_DATA_INTERLEAVE(HQM_SFI_RX_DATA_INTERLEAVE),
        .HQM_SFI_RX_DATA_LAYER_EN(HQM_SFI_RX_DATA_LAYER_EN),
        .HQM_SFI_RX_DATA_PARITY_EN(HQM_SFI_RX_DATA_PARITY_EN),
        .HQM_SFI_RX_DATA_PASS_HDR(HQM_SFI_RX_DATA_PASS_HDR),
        .HQM_SFI_RX_DATA_MAX_FC_VC(HQM_SFI_RX_DATA_MAX_FC_VC),
        .HQM_SFI_RX_DS(HQM_SFI_RX_DS),
        .HQM_SFI_RX_ECRC_SUPPORT(HQM_SFI_RX_ECRC_SUPPORT),
        .HQM_SFI_RX_FLIT_MODE_PREFIX_EN(HQM_SFI_RX_FLIT_MODE_PREFIX_EN),
        .HQM_SFI_RX_FATAL_EN(HQM_SFI_RX_FATAL_EN),
        .HQM_SFI_RX_H(HQM_SFI_RX_H),
        .HQM_SFI_RX_HDR_DATA_SEP(HQM_SFI_RX_HDR_DATA_SEP),
        .HQM_SFI_RX_HDR_MAX_FC_VC(HQM_SFI_RX_HDR_MAX_FC_VC),
        .HQM_SFI_RX_HGRAN(HQM_SFI_RX_HGRAN),
        .HQM_SFI_RX_HPARITY(HQM_SFI_RX_HPARITY),
        .HQM_SFI_RX_IDE_SUPPORT(HQM_SFI_RX_IDE_SUPPORT),
        .HQM_SFI_RX_M(HQM_SFI_RX_M),
        .HQM_SFI_RX_MAX_CRD_CNT_WIDTH(HQM_SFI_RX_MAX_CRD_CNT_WIDTH),
        .HQM_SFI_RX_MAX_HDR_WIDTH(HQM_SFI_RX_MAX_HDR_WIDTH),
        .HQM_SFI_RX_NDCRD(HQM_SFI_RX_NDCRD),
        .HQM_SFI_RX_NHCRD(HQM_SFI_RX_NHCRD),
        .HQM_SFI_RX_NUM_SHARED_POOLS(HQM_SFI_RX_NUM_SHARED_POOLS),
        .HQM_SFI_RX_PCIE_MERGED_SELECT(HQM_SFI_RX_PCIE_MERGED_SELECT),
        .HQM_SFI_RX_PCIE_SHARED_SELECT(HQM_SFI_RX_PCIE_SHARED_SELECT),
        .HQM_SFI_RX_RBN(HQM_SFI_RX_RBN),
        .HQM_SFI_RX_SH_DATA_CRD_BLK_SZ(HQM_SFI_RX_SH_DATA_CRD_BLK_SZ),
        .HQM_SFI_RX_SH_HDR_CRD_BLK_SZ(HQM_SFI_RX_SH_HDR_CRD_BLK_SZ),
        .HQM_SFI_RX_SHARED_CREDIT_EN(HQM_SFI_RX_SHARED_CREDIT_EN),
        .HQM_SFI_RX_TBN(HQM_SFI_RX_TBN),
        .HQM_SFI_RX_TX_CRD_REG(HQM_SFI_RX_TX_CRD_REG),
        .HQM_SFI_RX_VIRAL_EN(HQM_SFI_RX_VIRAL_EN),
        .HQM_SFI_RX_VR(HQM_SFI_RX_VR),
        .HQM_SFI_RX_VT(HQM_SFI_RX_VT),
        .HQM_SFI_TX_BCM_EN(HQM_SFI_TX_BCM_EN),
        .HQM_SFI_TX_BLOCK_EARLY_VLD_EN(HQM_SFI_TX_BLOCK_EARLY_VLD_EN),
        .HQM_SFI_TX_D(HQM_SFI_TX_D),
        .HQM_SFI_TX_DATA_AUX_PARITY_EN(HQM_SFI_TX_DATA_AUX_PARITY_EN),
        .HQM_SFI_TX_DATA_CRD_GRAN(HQM_SFI_TX_DATA_CRD_GRAN),
        .HQM_SFI_TX_DATA_INTERLEAVE(HQM_SFI_TX_DATA_INTERLEAVE),
        .HQM_SFI_TX_DATA_LAYER_EN(HQM_SFI_TX_DATA_LAYER_EN),
        .HQM_SFI_TX_DATA_PARITY_EN(HQM_SFI_TX_DATA_PARITY_EN),
        .HQM_SFI_TX_DATA_PASS_HDR(HQM_SFI_TX_DATA_PASS_HDR),
        .HQM_SFI_TX_DATA_MAX_FC_VC(HQM_SFI_TX_DATA_MAX_FC_VC),
        .HQM_SFI_TX_DS(HQM_SFI_TX_DS),
        .HQM_SFI_TX_ECRC_SUPPORT(HQM_SFI_TX_ECRC_SUPPORT),
        .HQM_SFI_TX_FLIT_MODE_PREFIX_EN(HQM_SFI_TX_FLIT_MODE_PREFIX_EN),
        .HQM_SFI_TX_FATAL_EN(HQM_SFI_TX_FATAL_EN),
        .HQM_SFI_TX_H(HQM_SFI_TX_H),
        .HQM_SFI_TX_HDR_DATA_SEP(HQM_SFI_TX_HDR_DATA_SEP),
        .HQM_SFI_TX_HDR_MAX_FC_VC(HQM_SFI_TX_HDR_MAX_FC_VC),
        .HQM_SFI_TX_HGRAN(HQM_SFI_TX_HGRAN),
        .HQM_SFI_TX_HPARITY(HQM_SFI_TX_HPARITY),
        .HQM_SFI_TX_IDE_SUPPORT(HQM_SFI_TX_IDE_SUPPORT),
        .HQM_SFI_TX_M(HQM_SFI_TX_M),
        .HQM_SFI_TX_MAX_CRD_CNT_WIDTH(HQM_SFI_TX_MAX_CRD_CNT_WIDTH),
        .HQM_SFI_TX_MAX_HDR_WIDTH(HQM_SFI_TX_MAX_HDR_WIDTH),
        .HQM_SFI_TX_NDCRD(HQM_SFI_TX_NDCRD),
        .HQM_SFI_TX_NHCRD(HQM_SFI_TX_NHCRD),
        .HQM_SFI_TX_NUM_SHARED_POOLS(HQM_SFI_TX_NUM_SHARED_POOLS),
        .HQM_SFI_TX_PCIE_MERGED_SELECT(HQM_SFI_TX_PCIE_MERGED_SELECT),
        .HQM_SFI_TX_PCIE_SHARED_SELECT(HQM_SFI_TX_PCIE_SHARED_SELECT),
        .HQM_SFI_TX_RBN(HQM_SFI_TX_RBN),
        .HQM_SFI_TX_SH_DATA_CRD_BLK_SZ(HQM_SFI_TX_SH_DATA_CRD_BLK_SZ),
        .HQM_SFI_TX_SH_HDR_CRD_BLK_SZ(HQM_SFI_TX_SH_HDR_CRD_BLK_SZ),
        .HQM_SFI_TX_SHARED_CREDIT_EN(HQM_SFI_TX_SHARED_CREDIT_EN),
        .HQM_SFI_TX_TBN(HQM_SFI_TX_TBN),
        .HQM_SFI_TX_TX_CRD_REG(HQM_SFI_TX_TX_CRD_REG),
        .HQM_SFI_TX_VIRAL_EN(HQM_SFI_TX_VIRAL_EN),
        .HQM_SFI_TX_VR(HQM_SFI_TX_VR),
        .HQM_SFI_TX_VT(HQM_SFI_TX_VT)) i_hqm_sif
      (.pgcb_clk                         (iosf_pgcb_clk),
       .powergood_rst_b,
       .pma_safemode,
       .hqm_inp_gated_clk,
       .hqm_gated_rst_b                  (hqm_gated_rst_b_mstr),
       // Tie to constant value: zero
       .strap_hqm_is_reg_ep              (1'b0),
       .strap_hqm_csr_cp,
       .strap_hqm_csr_rac,
       .strap_hqm_csr_wac,
       .strap_hqm_device_id,
       .strap_hqm_err_sb_dstid,
       .strap_hqm_err_sb_sai,
       .strap_hqm_tx_sai,
       .strap_hqm_cmpl_sai,
       .strap_hqm_resetprep_ack_sai,
       .strap_hqm_resetprep_sai_0,
       .strap_hqm_resetprep_sai_1,
       .strap_hqm_force_pok_sai_0,
       .strap_hqm_force_pok_sai_1,
       .strap_hqm_gpsb_srcid,
       .strap_hqm_16b_portids,
       .strap_hqm_do_serr_dstid,
       .strap_hqm_do_serr_tag,
       .strap_hqm_do_serr_sairs_valid,
       .strap_hqm_do_serr_sai,
       .strap_hqm_do_serr_rs,
       .side_pok,
       .side_clk,
       .side_clkreq,
       .side_clkack,
       .side_rst_b,
       .gpsb_side_ism_fabric,
       .gpsb_side_ism_agent,
       .side_pwrgate_pmc_wake,
       .gpsb_mpccup,
       .gpsb_mnpcup,
       .gpsb_mpcput,
       .gpsb_mnpput,
       .gpsb_meom,
       .gpsb_mpayload,
       .gpsb_mparity,
       .gpsb_tpccup,
       .gpsb_tnpcup,
       .gpsb_tpcput,
       .gpsb_tnpput,
       .gpsb_teom,
       .gpsb_tpayload,
       .gpsb_tparity,
       .sfi_tx_txcon_req,
       .sfi_tx_rxcon_ack,
       .sfi_tx_rxdiscon_nack,
       .sfi_tx_rx_empty,
       .sfi_tx_hdr_valid,
       .sfi_tx_hdr_early_valid,
       .sfi_tx_hdr_info_bytes,
       .sfi_tx_header,
       .sfi_tx_hdr_block,
       .sfi_tx_hdr_crd_rtn_valid,
       .sfi_tx_hdr_crd_rtn_vc_id,
       .sfi_tx_hdr_crd_rtn_fc_id,
       .sfi_tx_hdr_crd_rtn_value,
       .sfi_tx_hdr_crd_rtn_block,
       .sfi_tx_data_valid,
       .sfi_tx_data_early_valid,
       .sfi_tx_data_aux_parity,
       .sfi_tx_data_parity,
       .sfi_tx_data_poison,
       .sfi_tx_data_edb,
       .sfi_tx_data_start,
       .sfi_tx_data_end,
       .sfi_tx_data_info_byte,
       .sfi_tx_data,
       .sfi_tx_data_block,
       .sfi_tx_data_crd_rtn_valid,
       .sfi_tx_data_crd_rtn_vc_id,
       .sfi_tx_data_crd_rtn_fc_id,
       .sfi_tx_data_crd_rtn_value,
       .sfi_tx_data_crd_rtn_block,
       .sfi_rx_txcon_req,
       .sfi_rx_rxcon_ack,
       .sfi_rx_rxdiscon_nack,
       .sfi_rx_rx_empty,
       .sfi_rx_hdr_valid,
       .sfi_rx_hdr_early_valid,
       .sfi_rx_hdr_info_bytes,
       .sfi_rx_header,
       .sfi_rx_hdr_block,
       .sfi_rx_hdr_crd_rtn_valid,
       .sfi_rx_hdr_crd_rtn_vc_id,
       .sfi_rx_hdr_crd_rtn_fc_id,
       .sfi_rx_hdr_crd_rtn_value,
       .sfi_rx_hdr_crd_rtn_block,
       .sfi_rx_data_valid,
       .sfi_rx_data_early_valid,
       .sfi_rx_data_aux_parity,
       .sfi_rx_data_parity,
       .sfi_rx_data_poison,
       .sfi_rx_data_edb,
       .sfi_rx_data_start,
       .sfi_rx_data_end,
       .sfi_rx_data_info_byte,
       .sfi_rx_data,
       .sfi_rx_data_block,
       .sfi_rx_data_crd_rtn_valid,
       .sfi_rx_data_crd_rtn_vc_id,
       .sfi_rx_data_crd_rtn_fc_id,
       .sfi_rx_data_crd_rtn_value,
       .sfi_rx_data_crd_rtn_block,
       .prim_pwrgate_pmc_wake,
       .prim_freerun_clk                 (prim_clk),
       .prim_gated_clk,
       .prim_nonflr_clk,
       .prim_clkack,
       .prim_clkreq,
       .prim_clk_enable                  (i_hqm_sif_prim_clk_enable),
       .prim_clk_enable_cdc,
       .prim_clk_enable_sys,
       .prim_clk_ungate                  (i_hqm_sif_prim_clk_ungate),
       .prim_rst_b,
       .prim_gated_rst_b,
       .flr_triggered,
       .psel,
       .penable,
       .pwrite,
       .paddr,
       .pwdata,
       .puser,
       .pready,
       .pslverr,
       .prdata,
       .prdata_par,
       .hcw_enq_in_ready,
       .hcw_enq_in_v,
       .hcw_enq_in_data,
       .write_buffer_mstr_ready,
       .write_buffer_mstr_v,
       .write_buffer_mstr,
       .sif_alarm_ready,
       .sif_alarm_v,
       .sif_alarm_data,
       .pci_cfg_sciov_en,
       .pci_cfg_pmsixctl_msie,
       .pci_cfg_pmsixctl_fm,
       .pm_state,
       .pm_fsm_d0tod3_ok,
       .pm_fsm_d3tod0_ok,
       .pm_fsm_in_run,
       .pm_allow_ing_drop,
       .hqm_proc_reset_done,
       .hqm_proc_idle                    (hqm_proc_clkreq_b),
       .hqm_flr_prep                     (hqm_shields_up),
       .master_ctl_load,
       .master_ctl,
       .fdfx_sbparity_def,
       .fscan_byprst_b,
       .fscan_clkungate,
       .fscan_clkungate_syn,
       .fscan_latchclosed_b,
       .fscan_latchopen,
       .fscan_mode,
       .fscan_rstbypen,
       .fscan_shiften,
       .prim_jta_force_clkreq            (rtdr_func_po_iosfsb_ism[2]),
       .prim_jta_force_creditreq         (rtdr_func_po_iosfsb_ism[3]),
       .prim_jta_force_idle              (rtdr_func_po_iosfsb_ism[5]),
       .prim_jta_force_notidle           (rtdr_func_po_iosfsb_ism[4]),
       .gpsb_jta_clkgate_ovrd            (rtdr_func_po_iosfsb_ism[11]),
       .gpsb_jta_force_clkreq            (rtdr_func_po_iosfsb_ism[12]),
       .gpsb_jta_force_creditreq         (rtdr_func_po_iosfsb_ism[13]),
       .gpsb_jta_force_idle              (rtdr_func_po_iosfsb_ism[15]),
       .gpsb_jta_force_notidle           (rtdr_func_po_iosfsb_ism[14]),
       .cdc_prim_jta_force_clkreq        (rtdr_func_po_iosfsb_ism[2]),
       .cdc_prim_jta_clkgate_ovrd        (rtdr_func_po_iosfsb_ism[1]),
       .cdc_side_jta_force_clkreq        (rtdr_func_po_iosfsb_ism[12]),
       .cdc_side_jta_clkgate_ovrd        (rtdr_func_po_iosfsb_ism[0]),
       .fuse_force_on,
       .fuse_proc_disable,
       .early_fuses,
       .ip_ready,
       .strap_no_mgmt_acks,
       .reset_prep_ack,
       .pm_hqm_adr_assert,
       .hqm_pm_adr_ack,
       .hqm_triggers                     (hqm_triggers_in),
       .hqm_sif_visa,
       .rf_ibcpl_data_fifo_re            (i_hqm_sif_rf_ibcpl_data_fifo_re),
       .rf_ibcpl_data_fifo_rclk          (i_hqm_sif_rf_ibcpl_data_fifo_rclk),
       .rf_ibcpl_data_fifo_rclk_rst_n    (i_hqm_sif_rf_ibcpl_data_fifo_rclk_rst_n),
       .rf_ibcpl_data_fifo_raddr         (i_hqm_sif_rf_ibcpl_data_fifo_raddr),
       .rf_ibcpl_data_fifo_waddr         (i_hqm_sif_rf_ibcpl_data_fifo_waddr),
       .rf_ibcpl_data_fifo_we            (i_hqm_sif_rf_ibcpl_data_fifo_we),
       .rf_ibcpl_data_fifo_wclk          (i_hqm_sif_rf_ibcpl_data_fifo_wclk),
       .rf_ibcpl_data_fifo_wclk_rst_n    (i_hqm_sif_rf_ibcpl_data_fifo_wclk_rst_n),
       .rf_ibcpl_data_fifo_wdata         (i_hqm_sif_rf_ibcpl_data_fifo_wdata),
       .rf_ibcpl_data_fifo_rdata         (i_hqm_sif_rf_ibcpl_data_fifo_rdata),
       .rf_ibcpl_hdr_fifo_re             (i_hqm_sif_rf_ibcpl_hdr_fifo_re),
       .rf_ibcpl_hdr_fifo_rclk           (i_hqm_sif_rf_ibcpl_hdr_fifo_rclk),
       .rf_ibcpl_hdr_fifo_rclk_rst_n     (i_hqm_sif_rf_ibcpl_hdr_fifo_rclk_rst_n),
       .rf_ibcpl_hdr_fifo_raddr          (i_hqm_sif_rf_ibcpl_hdr_fifo_raddr),
       .rf_ibcpl_hdr_fifo_waddr          (i_hqm_sif_rf_ibcpl_hdr_fifo_waddr),
       .rf_ibcpl_hdr_fifo_we             (i_hqm_sif_rf_ibcpl_hdr_fifo_we),
       .rf_ibcpl_hdr_fifo_wclk           (i_hqm_sif_rf_ibcpl_hdr_fifo_wclk),
       .rf_ibcpl_hdr_fifo_wclk_rst_n     (i_hqm_sif_rf_ibcpl_hdr_fifo_wclk_rst_n),
       .rf_ibcpl_hdr_fifo_wdata          (i_hqm_sif_rf_ibcpl_hdr_fifo_wdata),
       .rf_ibcpl_hdr_fifo_rdata          (i_hqm_sif_rf_ibcpl_hdr_fifo_rdata),
       .rf_mstr_ll_data0_re              (i_hqm_sif_rf_mstr_ll_data0_re),
       .rf_mstr_ll_data0_rclk            (i_hqm_sif_rf_mstr_ll_data0_rclk),
       .rf_mstr_ll_data0_rclk_rst_n      (i_hqm_sif_rf_mstr_ll_data0_rclk_rst_n),
       .rf_mstr_ll_data0_raddr           (i_hqm_sif_rf_mstr_ll_data0_raddr),
       .rf_mstr_ll_data0_waddr           (i_hqm_sif_rf_mstr_ll_data0_waddr),
       .rf_mstr_ll_data0_we              (i_hqm_sif_rf_mstr_ll_data0_we),
       .rf_mstr_ll_data0_wclk            (i_hqm_sif_rf_mstr_ll_data0_wclk),
       .rf_mstr_ll_data0_wclk_rst_n      (i_hqm_sif_rf_mstr_ll_data0_wclk_rst_n),
       .rf_mstr_ll_data0_wdata           (i_hqm_sif_rf_mstr_ll_data0_wdata),
       .rf_mstr_ll_data0_rdata           (i_hqm_sif_rf_mstr_ll_data0_rdata),
       .rf_mstr_ll_data1_re              (i_hqm_sif_rf_mstr_ll_data1_re),
       .rf_mstr_ll_data1_rclk            (i_hqm_sif_rf_mstr_ll_data1_rclk),
       .rf_mstr_ll_data1_rclk_rst_n      (i_hqm_sif_rf_mstr_ll_data1_rclk_rst_n),
       .rf_mstr_ll_data1_raddr           (i_hqm_sif_rf_mstr_ll_data1_raddr),
       .rf_mstr_ll_data1_waddr           (i_hqm_sif_rf_mstr_ll_data1_waddr),
       .rf_mstr_ll_data1_we              (i_hqm_sif_rf_mstr_ll_data1_we),
       .rf_mstr_ll_data1_wclk            (i_hqm_sif_rf_mstr_ll_data1_wclk),
       .rf_mstr_ll_data1_wclk_rst_n      (i_hqm_sif_rf_mstr_ll_data1_wclk_rst_n),
       .rf_mstr_ll_data1_wdata           (i_hqm_sif_rf_mstr_ll_data1_wdata),
       .rf_mstr_ll_data1_rdata           (i_hqm_sif_rf_mstr_ll_data1_rdata),
       .rf_mstr_ll_data2_re              (i_hqm_sif_rf_mstr_ll_data2_re),
       .rf_mstr_ll_data2_rclk            (i_hqm_sif_rf_mstr_ll_data2_rclk),
       .rf_mstr_ll_data2_rclk_rst_n      (i_hqm_sif_rf_mstr_ll_data2_rclk_rst_n),
       .rf_mstr_ll_data2_raddr           (i_hqm_sif_rf_mstr_ll_data2_raddr),
       .rf_mstr_ll_data2_waddr           (i_hqm_sif_rf_mstr_ll_data2_waddr),
       .rf_mstr_ll_data2_we              (i_hqm_sif_rf_mstr_ll_data2_we),
       .rf_mstr_ll_data2_wclk            (i_hqm_sif_rf_mstr_ll_data2_wclk),
       .rf_mstr_ll_data2_wclk_rst_n      (i_hqm_sif_rf_mstr_ll_data2_wclk_rst_n),
       .rf_mstr_ll_data2_wdata           (i_hqm_sif_rf_mstr_ll_data2_wdata),
       .rf_mstr_ll_data2_rdata           (i_hqm_sif_rf_mstr_ll_data2_rdata),
       .rf_mstr_ll_data3_re              (i_hqm_sif_rf_mstr_ll_data3_re),
       .rf_mstr_ll_data3_rclk            (i_hqm_sif_rf_mstr_ll_data3_rclk),
       .rf_mstr_ll_data3_rclk_rst_n      (i_hqm_sif_rf_mstr_ll_data3_rclk_rst_n),
       .rf_mstr_ll_data3_raddr           (i_hqm_sif_rf_mstr_ll_data3_raddr),
       .rf_mstr_ll_data3_waddr           (i_hqm_sif_rf_mstr_ll_data3_waddr),
       .rf_mstr_ll_data3_we              (i_hqm_sif_rf_mstr_ll_data3_we),
       .rf_mstr_ll_data3_wclk            (i_hqm_sif_rf_mstr_ll_data3_wclk),
       .rf_mstr_ll_data3_wclk_rst_n      (i_hqm_sif_rf_mstr_ll_data3_wclk_rst_n),
       .rf_mstr_ll_data3_wdata           (i_hqm_sif_rf_mstr_ll_data3_wdata),
       .rf_mstr_ll_data3_rdata           (i_hqm_sif_rf_mstr_ll_data3_rdata),
       .rf_mstr_ll_hdr_re                (i_hqm_sif_rf_mstr_ll_hdr_re),
       .rf_mstr_ll_hdr_rclk              (i_hqm_sif_rf_mstr_ll_hdr_rclk),
       .rf_mstr_ll_hdr_rclk_rst_n        (i_hqm_sif_rf_mstr_ll_hdr_rclk_rst_n),
       .rf_mstr_ll_hdr_raddr             (i_hqm_sif_rf_mstr_ll_hdr_raddr),
       .rf_mstr_ll_hdr_waddr             (i_hqm_sif_rf_mstr_ll_hdr_waddr),
       .rf_mstr_ll_hdr_we                (i_hqm_sif_rf_mstr_ll_hdr_we),
       .rf_mstr_ll_hdr_wclk              (i_hqm_sif_rf_mstr_ll_hdr_wclk),
       .rf_mstr_ll_hdr_wclk_rst_n        (i_hqm_sif_rf_mstr_ll_hdr_wclk_rst_n),
       .rf_mstr_ll_hdr_wdata             (i_hqm_sif_rf_mstr_ll_hdr_wdata),
       .rf_mstr_ll_hdr_rdata             (i_hqm_sif_rf_mstr_ll_hdr_rdata),
       .rf_mstr_ll_hpa_re                (i_hqm_sif_rf_mstr_ll_hpa_re),
       .rf_mstr_ll_hpa_rclk              (i_hqm_sif_rf_mstr_ll_hpa_rclk),
       .rf_mstr_ll_hpa_rclk_rst_n        (i_hqm_sif_rf_mstr_ll_hpa_rclk_rst_n),
       .rf_mstr_ll_hpa_raddr             (i_hqm_sif_rf_mstr_ll_hpa_raddr),
       .rf_mstr_ll_hpa_waddr             (i_hqm_sif_rf_mstr_ll_hpa_waddr),
       .rf_mstr_ll_hpa_we                (i_hqm_sif_rf_mstr_ll_hpa_we),
       .rf_mstr_ll_hpa_wclk              (i_hqm_sif_rf_mstr_ll_hpa_wclk),
       .rf_mstr_ll_hpa_wclk_rst_n        (i_hqm_sif_rf_mstr_ll_hpa_wclk_rst_n),
       .rf_mstr_ll_hpa_wdata             (i_hqm_sif_rf_mstr_ll_hpa_wdata),
       .rf_mstr_ll_hpa_rdata             (i_hqm_sif_rf_mstr_ll_hpa_rdata),
       .rf_ri_tlq_fifo_npdata_re         (i_hqm_sif_rf_ri_tlq_fifo_npdata_re),
       .rf_ri_tlq_fifo_npdata_rclk       (i_hqm_sif_rf_ri_tlq_fifo_npdata_rclk),
       .rf_ri_tlq_fifo_npdata_rclk_rst_n (i_hqm_sif_rf_ri_tlq_fifo_npdata_rclk_rst_n),
       .rf_ri_tlq_fifo_npdata_raddr      (i_hqm_sif_rf_ri_tlq_fifo_npdata_raddr),
       .rf_ri_tlq_fifo_npdata_waddr      (i_hqm_sif_rf_ri_tlq_fifo_npdata_waddr),
       .rf_ri_tlq_fifo_npdata_we         (i_hqm_sif_rf_ri_tlq_fifo_npdata_we),
       .rf_ri_tlq_fifo_npdata_wclk       (i_hqm_sif_rf_ri_tlq_fifo_npdata_wclk),
       .rf_ri_tlq_fifo_npdata_wclk_rst_n (i_hqm_sif_rf_ri_tlq_fifo_npdata_wclk_rst_n),
       .rf_ri_tlq_fifo_npdata_wdata      (i_hqm_sif_rf_ri_tlq_fifo_npdata_wdata),
       .rf_ri_tlq_fifo_npdata_rdata      (i_hqm_sif_rf_ri_tlq_fifo_npdata_rdata),
       .rf_ri_tlq_fifo_nphdr_re          (i_hqm_sif_rf_ri_tlq_fifo_nphdr_re),
       .rf_ri_tlq_fifo_nphdr_rclk        (i_hqm_sif_rf_ri_tlq_fifo_nphdr_rclk),
       .rf_ri_tlq_fifo_nphdr_rclk_rst_n  (i_hqm_sif_rf_ri_tlq_fifo_nphdr_rclk_rst_n),
       .rf_ri_tlq_fifo_nphdr_raddr       (i_hqm_sif_rf_ri_tlq_fifo_nphdr_raddr),
       .rf_ri_tlq_fifo_nphdr_waddr       (i_hqm_sif_rf_ri_tlq_fifo_nphdr_waddr),
       .rf_ri_tlq_fifo_nphdr_we          (i_hqm_sif_rf_ri_tlq_fifo_nphdr_we),
       .rf_ri_tlq_fifo_nphdr_wclk        (i_hqm_sif_rf_ri_tlq_fifo_nphdr_wclk),
       .rf_ri_tlq_fifo_nphdr_wclk_rst_n  (i_hqm_sif_rf_ri_tlq_fifo_nphdr_wclk_rst_n),
       .rf_ri_tlq_fifo_nphdr_wdata       (i_hqm_sif_rf_ri_tlq_fifo_nphdr_wdata),
       .rf_ri_tlq_fifo_nphdr_rdata       (i_hqm_sif_rf_ri_tlq_fifo_nphdr_rdata),
       .rf_ri_tlq_fifo_pdata_re          (i_hqm_sif_rf_ri_tlq_fifo_pdata_re),
       .rf_ri_tlq_fifo_pdata_rclk        (i_hqm_sif_rf_ri_tlq_fifo_pdata_rclk),
       .rf_ri_tlq_fifo_pdata_rclk_rst_n  (i_hqm_sif_rf_ri_tlq_fifo_pdata_rclk_rst_n),
       .rf_ri_tlq_fifo_pdata_raddr       (i_hqm_sif_rf_ri_tlq_fifo_pdata_raddr),
       .rf_ri_tlq_fifo_pdata_waddr       (i_hqm_sif_rf_ri_tlq_fifo_pdata_waddr),
       .rf_ri_tlq_fifo_pdata_we          (i_hqm_sif_rf_ri_tlq_fifo_pdata_we),
       .rf_ri_tlq_fifo_pdata_wclk        (i_hqm_sif_rf_ri_tlq_fifo_pdata_wclk),
       .rf_ri_tlq_fifo_pdata_wclk_rst_n  (i_hqm_sif_rf_ri_tlq_fifo_pdata_wclk_rst_n),
       .rf_ri_tlq_fifo_pdata_wdata       (i_hqm_sif_rf_ri_tlq_fifo_pdata_wdata),
       .rf_ri_tlq_fifo_pdata_rdata       (i_hqm_sif_rf_ri_tlq_fifo_pdata_rdata),
       .rf_ri_tlq_fifo_phdr_re           (i_hqm_sif_rf_ri_tlq_fifo_phdr_re),
       .rf_ri_tlq_fifo_phdr_rclk         (i_hqm_sif_rf_ri_tlq_fifo_phdr_rclk),
       .rf_ri_tlq_fifo_phdr_rclk_rst_n   (i_hqm_sif_rf_ri_tlq_fifo_phdr_rclk_rst_n),
       .rf_ri_tlq_fifo_phdr_raddr        (i_hqm_sif_rf_ri_tlq_fifo_phdr_raddr),
       .rf_ri_tlq_fifo_phdr_waddr        (i_hqm_sif_rf_ri_tlq_fifo_phdr_waddr),
       .rf_ri_tlq_fifo_phdr_we           (i_hqm_sif_rf_ri_tlq_fifo_phdr_we),
       .rf_ri_tlq_fifo_phdr_wclk         (i_hqm_sif_rf_ri_tlq_fifo_phdr_wclk),
       .rf_ri_tlq_fifo_phdr_wclk_rst_n   (i_hqm_sif_rf_ri_tlq_fifo_phdr_wclk_rst_n),
       .rf_ri_tlq_fifo_phdr_wdata        (i_hqm_sif_rf_ri_tlq_fifo_phdr_wdata),
       .rf_ri_tlq_fifo_phdr_rdata        (i_hqm_sif_rf_ri_tlq_fifo_phdr_rdata),
       .rf_scrbd_mem_re                  (i_hqm_sif_rf_scrbd_mem_re),
       .rf_scrbd_mem_rclk                (i_hqm_sif_rf_scrbd_mem_rclk),
       .rf_scrbd_mem_rclk_rst_n          (i_hqm_sif_rf_scrbd_mem_rclk_rst_n),
       .rf_scrbd_mem_raddr               (i_hqm_sif_rf_scrbd_mem_raddr),
       .rf_scrbd_mem_waddr               (i_hqm_sif_rf_scrbd_mem_waddr),
       .rf_scrbd_mem_we                  (i_hqm_sif_rf_scrbd_mem_we),
       .rf_scrbd_mem_wclk                (i_hqm_sif_rf_scrbd_mem_wclk),
       .rf_scrbd_mem_wclk_rst_n          (i_hqm_sif_rf_scrbd_mem_wclk_rst_n),
       .rf_scrbd_mem_wdata               (i_hqm_sif_rf_scrbd_mem_wdata),
       .rf_scrbd_mem_rdata               (i_hqm_sif_rf_scrbd_mem_rdata),
       .rf_tlb_data0_4k_re               (i_hqm_sif_rf_tlb_data0_4k_re),
       .rf_tlb_data0_4k_rclk             (i_hqm_sif_rf_tlb_data0_4k_rclk),
       .rf_tlb_data0_4k_rclk_rst_n       (i_hqm_sif_rf_tlb_data0_4k_rclk_rst_n),
       .rf_tlb_data0_4k_raddr            (i_hqm_sif_rf_tlb_data0_4k_raddr),
       .rf_tlb_data0_4k_waddr            (i_hqm_sif_rf_tlb_data0_4k_waddr),
       .rf_tlb_data0_4k_we               (i_hqm_sif_rf_tlb_data0_4k_we),
       .rf_tlb_data0_4k_wclk             (i_hqm_sif_rf_tlb_data0_4k_wclk),
       .rf_tlb_data0_4k_wclk_rst_n       (i_hqm_sif_rf_tlb_data0_4k_wclk_rst_n),
       .rf_tlb_data0_4k_wdata            (i_hqm_sif_rf_tlb_data0_4k_wdata),
       .rf_tlb_data0_4k_rdata            (i_hqm_sif_rf_tlb_data0_4k_rdata),
       .rf_tlb_data1_4k_re               (i_hqm_sif_rf_tlb_data1_4k_re),
       .rf_tlb_data1_4k_rclk             (i_hqm_sif_rf_tlb_data1_4k_rclk),
       .rf_tlb_data1_4k_rclk_rst_n       (i_hqm_sif_rf_tlb_data1_4k_rclk_rst_n),
       .rf_tlb_data1_4k_raddr            (i_hqm_sif_rf_tlb_data1_4k_raddr),
       .rf_tlb_data1_4k_waddr            (i_hqm_sif_rf_tlb_data1_4k_waddr),
       .rf_tlb_data1_4k_we               (i_hqm_sif_rf_tlb_data1_4k_we),
       .rf_tlb_data1_4k_wclk             (i_hqm_sif_rf_tlb_data1_4k_wclk),
       .rf_tlb_data1_4k_wclk_rst_n       (i_hqm_sif_rf_tlb_data1_4k_wclk_rst_n),
       .rf_tlb_data1_4k_wdata            (i_hqm_sif_rf_tlb_data1_4k_wdata),
       .rf_tlb_data1_4k_rdata            (i_hqm_sif_rf_tlb_data1_4k_rdata),
       .rf_tlb_data2_4k_re               (i_hqm_sif_rf_tlb_data2_4k_re),
       .rf_tlb_data2_4k_rclk             (i_hqm_sif_rf_tlb_data2_4k_rclk),
       .rf_tlb_data2_4k_rclk_rst_n       (i_hqm_sif_rf_tlb_data2_4k_rclk_rst_n),
       .rf_tlb_data2_4k_raddr            (i_hqm_sif_rf_tlb_data2_4k_raddr),
       .rf_tlb_data2_4k_waddr            (i_hqm_sif_rf_tlb_data2_4k_waddr),
       .rf_tlb_data2_4k_we               (i_hqm_sif_rf_tlb_data2_4k_we),
       .rf_tlb_data2_4k_wclk             (i_hqm_sif_rf_tlb_data2_4k_wclk),
       .rf_tlb_data2_4k_wclk_rst_n       (i_hqm_sif_rf_tlb_data2_4k_wclk_rst_n),
       .rf_tlb_data2_4k_wdata            (i_hqm_sif_rf_tlb_data2_4k_wdata),
       .rf_tlb_data2_4k_rdata            (i_hqm_sif_rf_tlb_data2_4k_rdata),
       .rf_tlb_data3_4k_re               (i_hqm_sif_rf_tlb_data3_4k_re),
       .rf_tlb_data3_4k_rclk             (i_hqm_sif_rf_tlb_data3_4k_rclk),
       .rf_tlb_data3_4k_rclk_rst_n       (i_hqm_sif_rf_tlb_data3_4k_rclk_rst_n),
       .rf_tlb_data3_4k_raddr            (i_hqm_sif_rf_tlb_data3_4k_raddr),
       .rf_tlb_data3_4k_waddr            (i_hqm_sif_rf_tlb_data3_4k_waddr),
       .rf_tlb_data3_4k_we               (i_hqm_sif_rf_tlb_data3_4k_we),
       .rf_tlb_data3_4k_wclk             (i_hqm_sif_rf_tlb_data3_4k_wclk),
       .rf_tlb_data3_4k_wclk_rst_n       (i_hqm_sif_rf_tlb_data3_4k_wclk_rst_n),
       .rf_tlb_data3_4k_wdata            (i_hqm_sif_rf_tlb_data3_4k_wdata),
       .rf_tlb_data3_4k_rdata            (i_hqm_sif_rf_tlb_data3_4k_rdata),
       .rf_tlb_data4_4k_re               (i_hqm_sif_rf_tlb_data4_4k_re),
       .rf_tlb_data4_4k_rclk             (i_hqm_sif_rf_tlb_data4_4k_rclk),
       .rf_tlb_data4_4k_rclk_rst_n       (i_hqm_sif_rf_tlb_data4_4k_rclk_rst_n),
       .rf_tlb_data4_4k_raddr            (i_hqm_sif_rf_tlb_data4_4k_raddr),
       .rf_tlb_data4_4k_waddr            (i_hqm_sif_rf_tlb_data4_4k_waddr),
       .rf_tlb_data4_4k_we               (i_hqm_sif_rf_tlb_data4_4k_we),
       .rf_tlb_data4_4k_wclk             (i_hqm_sif_rf_tlb_data4_4k_wclk),
       .rf_tlb_data4_4k_wclk_rst_n       (i_hqm_sif_rf_tlb_data4_4k_wclk_rst_n),
       .rf_tlb_data4_4k_wdata            (i_hqm_sif_rf_tlb_data4_4k_wdata),
       .rf_tlb_data4_4k_rdata            (i_hqm_sif_rf_tlb_data4_4k_rdata),
       .rf_tlb_data5_4k_re               (i_hqm_sif_rf_tlb_data5_4k_re),
       .rf_tlb_data5_4k_rclk             (i_hqm_sif_rf_tlb_data5_4k_rclk),
       .rf_tlb_data5_4k_rclk_rst_n       (i_hqm_sif_rf_tlb_data5_4k_rclk_rst_n),
       .rf_tlb_data5_4k_raddr            (i_hqm_sif_rf_tlb_data5_4k_raddr),
       .rf_tlb_data5_4k_waddr            (i_hqm_sif_rf_tlb_data5_4k_waddr),
       .rf_tlb_data5_4k_we               (i_hqm_sif_rf_tlb_data5_4k_we),
       .rf_tlb_data5_4k_wclk             (i_hqm_sif_rf_tlb_data5_4k_wclk),
       .rf_tlb_data5_4k_wclk_rst_n       (i_hqm_sif_rf_tlb_data5_4k_wclk_rst_n),
       .rf_tlb_data5_4k_wdata            (i_hqm_sif_rf_tlb_data5_4k_wdata),
       .rf_tlb_data5_4k_rdata            (i_hqm_sif_rf_tlb_data5_4k_rdata),
       .rf_tlb_data6_4k_re               (i_hqm_sif_rf_tlb_data6_4k_re),
       .rf_tlb_data6_4k_rclk             (i_hqm_sif_rf_tlb_data6_4k_rclk),
       .rf_tlb_data6_4k_rclk_rst_n       (i_hqm_sif_rf_tlb_data6_4k_rclk_rst_n),
       .rf_tlb_data6_4k_raddr            (i_hqm_sif_rf_tlb_data6_4k_raddr),
       .rf_tlb_data6_4k_waddr            (i_hqm_sif_rf_tlb_data6_4k_waddr),
       .rf_tlb_data6_4k_we               (i_hqm_sif_rf_tlb_data6_4k_we),
       .rf_tlb_data6_4k_wclk             (i_hqm_sif_rf_tlb_data6_4k_wclk),
       .rf_tlb_data6_4k_wclk_rst_n       (i_hqm_sif_rf_tlb_data6_4k_wclk_rst_n),
       .rf_tlb_data6_4k_wdata            (i_hqm_sif_rf_tlb_data6_4k_wdata),
       .rf_tlb_data6_4k_rdata            (i_hqm_sif_rf_tlb_data6_4k_rdata),
       .rf_tlb_data7_4k_re               (i_hqm_sif_rf_tlb_data7_4k_re),
       .rf_tlb_data7_4k_rclk             (i_hqm_sif_rf_tlb_data7_4k_rclk),
       .rf_tlb_data7_4k_rclk_rst_n       (i_hqm_sif_rf_tlb_data7_4k_rclk_rst_n),
       .rf_tlb_data7_4k_raddr            (i_hqm_sif_rf_tlb_data7_4k_raddr),
       .rf_tlb_data7_4k_waddr            (i_hqm_sif_rf_tlb_data7_4k_waddr),
       .rf_tlb_data7_4k_we               (i_hqm_sif_rf_tlb_data7_4k_we),
       .rf_tlb_data7_4k_wclk             (i_hqm_sif_rf_tlb_data7_4k_wclk),
       .rf_tlb_data7_4k_wclk_rst_n       (i_hqm_sif_rf_tlb_data7_4k_wclk_rst_n),
       .rf_tlb_data7_4k_wdata            (i_hqm_sif_rf_tlb_data7_4k_wdata),
       .rf_tlb_data7_4k_rdata            (i_hqm_sif_rf_tlb_data7_4k_rdata),
       .rf_tlb_tag0_4k_re                (i_hqm_sif_rf_tlb_tag0_4k_re),
       .rf_tlb_tag0_4k_rclk              (i_hqm_sif_rf_tlb_tag0_4k_rclk),
       .rf_tlb_tag0_4k_rclk_rst_n        (i_hqm_sif_rf_tlb_tag0_4k_rclk_rst_n),
       .rf_tlb_tag0_4k_raddr             (i_hqm_sif_rf_tlb_tag0_4k_raddr),
       .rf_tlb_tag0_4k_waddr             (i_hqm_sif_rf_tlb_tag0_4k_waddr),
       .rf_tlb_tag0_4k_we                (i_hqm_sif_rf_tlb_tag0_4k_we),
       .rf_tlb_tag0_4k_wclk              (i_hqm_sif_rf_tlb_tag0_4k_wclk),
       .rf_tlb_tag0_4k_wclk_rst_n        (i_hqm_sif_rf_tlb_tag0_4k_wclk_rst_n),
       .rf_tlb_tag0_4k_wdata             (i_hqm_sif_rf_tlb_tag0_4k_wdata),
       .rf_tlb_tag0_4k_rdata             (i_hqm_sif_rf_tlb_tag0_4k_rdata),
       .rf_tlb_tag1_4k_re                (i_hqm_sif_rf_tlb_tag1_4k_re),
       .rf_tlb_tag1_4k_rclk              (i_hqm_sif_rf_tlb_tag1_4k_rclk),
       .rf_tlb_tag1_4k_rclk_rst_n        (i_hqm_sif_rf_tlb_tag1_4k_rclk_rst_n),
       .rf_tlb_tag1_4k_raddr             (i_hqm_sif_rf_tlb_tag1_4k_raddr),
       .rf_tlb_tag1_4k_waddr             (i_hqm_sif_rf_tlb_tag1_4k_waddr),
       .rf_tlb_tag1_4k_we                (i_hqm_sif_rf_tlb_tag1_4k_we),
       .rf_tlb_tag1_4k_wclk              (i_hqm_sif_rf_tlb_tag1_4k_wclk),
       .rf_tlb_tag1_4k_wclk_rst_n        (i_hqm_sif_rf_tlb_tag1_4k_wclk_rst_n),
       .rf_tlb_tag1_4k_wdata             (i_hqm_sif_rf_tlb_tag1_4k_wdata),
       .rf_tlb_tag1_4k_rdata             (i_hqm_sif_rf_tlb_tag1_4k_rdata),
       .rf_tlb_tag2_4k_re                (i_hqm_sif_rf_tlb_tag2_4k_re),
       .rf_tlb_tag2_4k_rclk              (i_hqm_sif_rf_tlb_tag2_4k_rclk),
       .rf_tlb_tag2_4k_rclk_rst_n        (i_hqm_sif_rf_tlb_tag2_4k_rclk_rst_n),
       .rf_tlb_tag2_4k_raddr             (i_hqm_sif_rf_tlb_tag2_4k_raddr),
       .rf_tlb_tag2_4k_waddr             (i_hqm_sif_rf_tlb_tag2_4k_waddr),
       .rf_tlb_tag2_4k_we                (i_hqm_sif_rf_tlb_tag2_4k_we),
       .rf_tlb_tag2_4k_wclk              (i_hqm_sif_rf_tlb_tag2_4k_wclk),
       .rf_tlb_tag2_4k_wclk_rst_n        (i_hqm_sif_rf_tlb_tag2_4k_wclk_rst_n),
       .rf_tlb_tag2_4k_wdata             (i_hqm_sif_rf_tlb_tag2_4k_wdata),
       .rf_tlb_tag2_4k_rdata             (i_hqm_sif_rf_tlb_tag2_4k_rdata),
       .rf_tlb_tag3_4k_re                (i_hqm_sif_rf_tlb_tag3_4k_re),
       .rf_tlb_tag3_4k_rclk              (i_hqm_sif_rf_tlb_tag3_4k_rclk),
       .rf_tlb_tag3_4k_rclk_rst_n        (i_hqm_sif_rf_tlb_tag3_4k_rclk_rst_n),
       .rf_tlb_tag3_4k_raddr             (i_hqm_sif_rf_tlb_tag3_4k_raddr),
       .rf_tlb_tag3_4k_waddr             (i_hqm_sif_rf_tlb_tag3_4k_waddr),
       .rf_tlb_tag3_4k_we                (i_hqm_sif_rf_tlb_tag3_4k_we),
       .rf_tlb_tag3_4k_wclk              (i_hqm_sif_rf_tlb_tag3_4k_wclk),
       .rf_tlb_tag3_4k_wclk_rst_n        (i_hqm_sif_rf_tlb_tag3_4k_wclk_rst_n),
       .rf_tlb_tag3_4k_wdata             (i_hqm_sif_rf_tlb_tag3_4k_wdata),
       .rf_tlb_tag3_4k_rdata             (i_hqm_sif_rf_tlb_tag3_4k_rdata),
       .rf_tlb_tag4_4k_re                (i_hqm_sif_rf_tlb_tag4_4k_re),
       .rf_tlb_tag4_4k_rclk              (i_hqm_sif_rf_tlb_tag4_4k_rclk),
       .rf_tlb_tag4_4k_rclk_rst_n        (i_hqm_sif_rf_tlb_tag4_4k_rclk_rst_n),
       .rf_tlb_tag4_4k_raddr             (i_hqm_sif_rf_tlb_tag4_4k_raddr),
       .rf_tlb_tag4_4k_waddr             (i_hqm_sif_rf_tlb_tag4_4k_waddr),
       .rf_tlb_tag4_4k_we                (i_hqm_sif_rf_tlb_tag4_4k_we),
       .rf_tlb_tag4_4k_wclk              (i_hqm_sif_rf_tlb_tag4_4k_wclk),
       .rf_tlb_tag4_4k_wclk_rst_n        (i_hqm_sif_rf_tlb_tag4_4k_wclk_rst_n),
       .rf_tlb_tag4_4k_wdata             (i_hqm_sif_rf_tlb_tag4_4k_wdata),
       .rf_tlb_tag4_4k_rdata             (i_hqm_sif_rf_tlb_tag4_4k_rdata),
       .rf_tlb_tag5_4k_re                (i_hqm_sif_rf_tlb_tag5_4k_re),
       .rf_tlb_tag5_4k_rclk              (i_hqm_sif_rf_tlb_tag5_4k_rclk),
       .rf_tlb_tag5_4k_rclk_rst_n        (i_hqm_sif_rf_tlb_tag5_4k_rclk_rst_n),
       .rf_tlb_tag5_4k_raddr             (i_hqm_sif_rf_tlb_tag5_4k_raddr),
       .rf_tlb_tag5_4k_waddr             (i_hqm_sif_rf_tlb_tag5_4k_waddr),
       .rf_tlb_tag5_4k_we                (i_hqm_sif_rf_tlb_tag5_4k_we),
       .rf_tlb_tag5_4k_wclk              (i_hqm_sif_rf_tlb_tag5_4k_wclk),
       .rf_tlb_tag5_4k_wclk_rst_n        (i_hqm_sif_rf_tlb_tag5_4k_wclk_rst_n),
       .rf_tlb_tag5_4k_wdata             (i_hqm_sif_rf_tlb_tag5_4k_wdata),
       .rf_tlb_tag5_4k_rdata             (i_hqm_sif_rf_tlb_tag5_4k_rdata),
       .rf_tlb_tag6_4k_re                (i_hqm_sif_rf_tlb_tag6_4k_re),
       .rf_tlb_tag6_4k_rclk              (i_hqm_sif_rf_tlb_tag6_4k_rclk),
       .rf_tlb_tag6_4k_rclk_rst_n        (i_hqm_sif_rf_tlb_tag6_4k_rclk_rst_n),
       .rf_tlb_tag6_4k_raddr             (i_hqm_sif_rf_tlb_tag6_4k_raddr),
       .rf_tlb_tag6_4k_waddr             (i_hqm_sif_rf_tlb_tag6_4k_waddr),
       .rf_tlb_tag6_4k_we                (i_hqm_sif_rf_tlb_tag6_4k_we),
       .rf_tlb_tag6_4k_wclk              (i_hqm_sif_rf_tlb_tag6_4k_wclk),
       .rf_tlb_tag6_4k_wclk_rst_n        (i_hqm_sif_rf_tlb_tag6_4k_wclk_rst_n),
       .rf_tlb_tag6_4k_wdata             (i_hqm_sif_rf_tlb_tag6_4k_wdata),
       .rf_tlb_tag6_4k_rdata             (i_hqm_sif_rf_tlb_tag6_4k_rdata),
       .rf_tlb_tag7_4k_re                (i_hqm_sif_rf_tlb_tag7_4k_re),
       .rf_tlb_tag7_4k_rclk              (i_hqm_sif_rf_tlb_tag7_4k_rclk),
       .rf_tlb_tag7_4k_rclk_rst_n        (i_hqm_sif_rf_tlb_tag7_4k_rclk_rst_n),
       .rf_tlb_tag7_4k_raddr             (i_hqm_sif_rf_tlb_tag7_4k_raddr),
       .rf_tlb_tag7_4k_waddr             (i_hqm_sif_rf_tlb_tag7_4k_waddr),
       .rf_tlb_tag7_4k_we                (i_hqm_sif_rf_tlb_tag7_4k_we),
       .rf_tlb_tag7_4k_wclk              (i_hqm_sif_rf_tlb_tag7_4k_wclk),
       .rf_tlb_tag7_4k_wclk_rst_n        (i_hqm_sif_rf_tlb_tag7_4k_wclk_rst_n),
       .rf_tlb_tag7_4k_wdata             (i_hqm_sif_rf_tlb_tag7_4k_wdata),
       .rf_tlb_tag7_4k_rdata             (i_hqm_sif_rf_tlb_tag7_4k_rdata));

   hqm_AW_flop i_hqm_sif_nonflr_clk_enable_rptr
      (.clk    (prim_clk),
       .rst_n  (side_rst_sync_prim_n),
       .data   (prim_clk_enable_cdc),
       .data_q (nonflr_clk_enable_rptr));

   hqm_AW_flop i_hqm_sif_prim_clk_enable_rptr
      (.clk    (prim_clk),
       .rst_n  (side_rst_sync_prim_n),
       .data   (prim_clk_enable_sys),
       .data_q (prim_clk_enable_rptr));

   hqm_AW_clkgate i_hqm_sif_prim_clkgate
      (.clk             (prim_clk),
       .enable          (prim_clk_enable_rptr),
       .cfg_clkungate   (prim_clk_ungate_rptr),
       .fscan_clkungate,
       .gated_clk       (prim_gated_clk));

   hqm_AW_clkgate i_hqm_sif_prim_clknonflr
      (.clk             (prim_clk),
       .enable          (nonflr_clk_enable_rptr),
       .cfg_clkungate   (prim_clk_ungate_rptr),
       .fscan_clkungate,
       .gated_clk       (prim_nonflr_clk));

   hqm_visa
      #(.HQM_DTF_TO_CNT_THRESHOLD(HQM_DTF_TO_CNT_THRESHOLD),
        .HQM_DTF_DATA_WIDTH(HQM_DTF_DATA_WIDTH),
        .HQM_TRIGFABWIDTH(HQM_TRIGFABWIDTH),
        .HQM_DVP_USE_PUSH_SWD(HQM_DVP_USE_PUSH_SWD),
        .HQM_DVP_USE_LEGACY_TIMESTAMP(HQM_DVP_USE_LEGACY_TIMESTAMP),
        .HQM_DTF_HEADER_WIDTH(HQM_DTF_HEADER_WIDTH)) i_hqm_visa
      (// Tie to constant value: 0
       .fvisa_frame_vcfn          (1'b0),
       // Tie to constant value: 0
       .fvisa_serdata_vcfn        (1'b0),
       // Tie to constant value: 0
       .fvisa_serstb_vcfn         (1'b0),
       // Tie to constant value: 0
       .fvisa_startid0_vcfn       (9'b0),
       // Tie to constant value: 0
       .fvisa_startid1_vcfn       (9'b0),
       // Tie to constant value: 0
       .fvisa_startid2_vcfn       (9'b0),
       // Tie to constant value: 0
       .fvisa_startid3_vcfn       (9'b0),
       .prim_freerun_clk          (prim_clk),
       .powergood_rst_b,
       // Tie to constant value: 0
       .visa_all_dis              (1'b0),
       // Tie to constant value: 0
       .visa_customer_dis         (1'b0),
       .avisa_dbgbus0_vcfn        (),
       .avisa_dbgbus1_vcfn        (),
       .avisa_dbgbus2_vcfn        (),
       .avisa_dbgbus3_vcfn        (),
       .hqm_sif_visa,
       .pgcb_clk,
       .hqm_cdc_visa,
       .hqm_pgcbunit_visa         (hqm_pgcb_visa),
       .hqm_pmsm_visa,
       .clk                       (i_system_buf_hqm_clk_trunk_o),
       .hqm_system_visa_str,
       .side_clk,
       .wd_clkreq,
       .hqm_cfg_master_clkreq_b   (i_hqm_master_hqm_cfg_master_clkreq_b),
       .side_rst_b,
       .prim_gated_rst_b,
       .hqm_gated_rst_b           (hqm_gated_rst_b_mstr),
       .hqm_clk_rptr_rst_b        (i_hqm_master_hqm_clk_rptr_rst_b),
       .hqm_pwrgood_rst_b         (hqm_pwrgood_rst_b_internal),
       .prochot,
       .master_ctl,
       .pgcb_isol_en_b,
       .pgcb_isol_en              (i_hqm_master_pgcb_isol_en),
       .pgcb_fet_en_b             (i_hqm_master_pgcb_fet_en_b),
       .pgcb_fet_en_ack_b,
       // Tie to constant value: 0
       .pgcb_fet_en_ack_b_sys     (1'b0),
       // Tie to constant value: 0
       .pgcb_fet_en_ack_b_qed     (1'b0),
       .cdc_hqm_jta_force_clkreq  (rtdr_func_po_iosfsb_ism[2]),
       .cdc_hqm_jta_clkgate_ovrd  (rtdr_func_po_iosfsb_ism[1]),
       .hqm_fullrate_clk          (i_system_buf_hqm_clk_trunk_o),
       // Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: one
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  dqed_cfg_req_down_read
       //  dqed_cfg_req_down_write
       //  dqed_cfg_req_down
       //  dqed_cfg_rsp_down_ack
       //  dqed_cfg_rsp_down
       //  Tie to constant value: zero
       //  Tie to constant value: zero
       //  qed_alarm_down_v
       //  qed_alarm_down_ready
       //  dqed_alarm_down_v
       //  dqed_alarm_down_ready
       .hqm_core_visa_str         ({ap_alarm_up_ready, 
                                    aqed_alarm_down_v, 
                                    4'b0, 
                                    i_hqm_visa_hqm_core_visa_str_253, 
                                    i_hqm_visa_hqm_core_visa_str_252, 
                                    lsp_alarm_up_ready, 
                                    ap_alarm_down_v, 
                                    rop_alarm_up_ready, 
                                    qed_alarm_down_v, 
                                    qed_alarm_up_ready, 
                                    lsp_alarm_down_v, 
                                    chp_alarm_up_ready, 
                                    rop_alarm_down_v, 
                                    2'b0, 
                                    i_hqm_visa_hqm_core_visa_str_241_240[1:0], 
                                    aqed_cfg_rsp_down_ack, 
                                    i_hqm_visa_hqm_core_visa_str_238_237[1:0], 
                                    aqed_cfg_req_down_write, 
                                    aqed_cfg_req_down_read, 
                                    7'b0, 
                                    i_hqm_visa_hqm_core_visa_str_227_226[1:0], 
                                    qed_cfg_rsp_down_ack, 
                                    i_hqm_visa_hqm_core_visa_str_224_223[1:0], 
                                    qed_cfg_req_down_write, 
                                    qed_cfg_req_down_read, 
                                    7'b0, 
                                    i_hqm_visa_hqm_core_visa_str_213_212[1:0], 
                                    ap_cfg_rsp_down_ack, 
                                    i_hqm_visa_hqm_core_visa_str_210_209[1:0], 
                                    ap_cfg_req_down_write, 
                                    ap_cfg_req_down_read, 
                                    7'b0, 
                                    i_hqm_visa_hqm_core_visa_str_199_198[1:0], 
                                    lsp_cfg_rsp_down_ack, 
                                    i_hqm_visa_hqm_core_visa_str_196_195[1:0], 
                                    lsp_cfg_req_down_write, 
                                    lsp_cfg_req_down_read, 
                                    i_hqm_visa_hqm_core_visa_str_192_191[1:0], 
                                    rop_cfg_rsp_down_ack, 
                                    i_hqm_visa_hqm_core_visa_str_189_188[1:0], 
                                    rop_cfg_req_down_write, 
                                    rop_cfg_req_down_read, 
                                    i_hqm_visa_hqm_core_visa_str_185_184[1:0], 
                                    chp_cfg_rsp_down_ack, 
                                    i_hqm_visa_hqm_core_visa_str_182_181[1:0], 
                                    chp_cfg_req_down_write, 
                                    chp_cfg_req_down_read, 
                                    i_hqm_visa_hqm_core_visa_str_178_177[1:0], 
                                    system_cfg_rsp_down_ack, 
                                    i_hqm_visa_hqm_core_visa_str_175_174[1:0], 
                                    system_cfg_req_down_write, 
                                    system_cfg_req_down_read, 
                                    rop_lsp_reordercmp_ready, 
                                    rop_lsp_reordercmp_v, 
                                    aqed_lsp_sch_ready, 
                                    aqed_lsp_sch_v, 
                                    aqed_chp_sch_ready, 
                                    aqed_chp_sch_v, 
                                    aqed_ap_enq_ready, 
                                    aqed_ap_enq_v, 
                                    2'b0, 
                                    qed_aqed_enq_ready, 
                                    qed_aqed_enq_v, 
                                    qed_chp_sch_ready, 
                                    qed_chp_sch_v, 
                                    ap_aqed_ready, 
                                    ap_aqed_v, 
                                    2'b0, 
                                    dp_lsp_enq_rorply_ready, 
                                    dp_lsp_enq_rorply_v, 
                                    dp_lsp_enq_dir_ready, 
                                    dp_lsp_enq_dir_v, 
                                    2'b0, 
                                    nalb_lsp_enq_rorply_ready, 
                                    nalb_lsp_enq_rorply_v, 
                                    nalb_lsp_enq_lb_ready, 
                                    nalb_lsp_enq_lb_v, 
                                    lsp_nalb_sch_atq_ready, 
                                    lsp_nalb_sch_atq_v, 
                                    lsp_dp_sch_rorply_ready, 
                                    lsp_dp_sch_rorply_v, 
                                    lsp_nalb_sch_rorply_ready, 
                                    lsp_nalb_sch_rorply_v, 
                                    lsp_dp_sch_dir_ready, 
                                    lsp_dp_sch_dir_v, 
                                    lsp_nalb_sch_unoord_ready, 
                                    lsp_nalb_sch_unoord_v, 
                                    rop_dqed_enq_ready, 
                                    rop_qed_enq_ready, 
                                    rop_qed_dqed_enq_v, 
                                    rop_nalb_enq_ready, 
                                    rop_nalb_enq_v, 
                                    rop_dp_enq_ready, 
                                    rop_dp_enq_v, 
                                    chp_lsp_token_ready, 
                                    chp_lsp_token_v, 
                                    visa_str_chp_lsp_cmp_data, 
                                    chp_lsp_cmp_ready, 
                                    chp_lsp_cmp_v, 
                                    chp_rop_hcw_ready, 
                                    chp_rop_hcw_v, 
                                    6'b0, 
                                    hcw_sched_w_req_ready, 
                                    hcw_sched_w_req_valid, 
                                    4'b0, 
                                    hcw_enq_w_req_ready, 
                                    hcw_enq_w_req_valid, 
                                    2'b0, 
                                    cwdi_interrupt_w_req_ready, 
                                    cwdi_interrupt_w_req_valid, 
                                    interrupt_w_req_ready, 
                                    interrupt_w_req_valid, 
                                    1'b0, 
                                    aqed_unit_pipeidle, 
                                    qed_unit_pipeidle, 
                                    dp_unit_pipeidle, 
                                    ap_unit_pipeidle, 
                                    nalb_unit_pipeidle, 
                                    lsp_unit_pipeidle, 
                                    rop_unit_pipeidle, 
                                    chp_unit_pipeidle, 
                                    system_idle, 
                                    aqed_unit_idle, 
                                    qed_unit_idle, 
                                    dp_unit_idle, 
                                    ap_unit_idle, 
                                    nalb_unit_idle, 
                                    lsp_unit_idle, 
                                    rop_unit_idle, 
                                    chp_unit_idle, 
                                    3'b0, 
                                    hqm_proc_clk_en_sys, 
                                    hqm_proc_clk_en_nalb, 
                                    hqm_proc_clk_en_dir, 
                                    hqm_proc_clk_en_qed, 
                                    hqm_proc_clk_en_lsp, 
                                    hqm_proc_clk_en_chp, 
                                    system_reset_done, 
                                    aqed_reset_done, 
                                    qed_reset_done, 
                                    dp_reset_done, 
                                    ap_reset_done, 
                                    nalb_reset_done, 
                                    lsp_reset_done, 
                                    rop_reset_done, 
                                    chp_reset_done, 
                                    15'b0, 
                                    hqm_alarm_v, 
                                    hqm_alarm_ready, 
                                    visa_str_hqm_proc_pipeidle, 
                                    visa_str_hqm_proc_idle, 
                                    1'b1, 
                                    rop_qed_force_clockon, 
                                    i_hqm_master_hqm_proc_reset_done_sync_hqm, 
                                    26'b0, 
                                    visa_str_pm_ip_clk_halt_b_2_rpt_0_iosf, 
                                    visa_str_hqm_flr_prep, 
                                    visa_str_hqm_gated_local_override, 
                                    visa_str_hqm_cdc_clk_enable, 
                                    visa_str_hqm_gclock_enable, 
                                    visa_str_hqm_clk_throttle, 
                                    visa_str_hqm_clk_enable, 
                                    visa_str_prim_clk_enable, 
                                    7'b0, 
                                    hqm_gated_rst_b_mstr}),
       .fscan_byprst_b,
       .fscan_rstbypen,
       .fscan_mode,
       .fdtf_clk,
       .fdtf_cry_clk,
       .fdtf_rst_b,
       .pma_safemode,
       .fdtf_survive_mode,
       .fdtf_fast_cnt_width,
       .fdtf_packetizer_mid,
       .fdtf_packetizer_cid,
       .adtf_dnstream_header,
       .adtf_dnstream_data,
       .adtf_dnstream_valid,
       .fdtf_upstream_credit,
       .fdtf_upstream_active,
       .fdtf_upstream_sync,
       .fdtf_serial_download_tsc,
       .fdtf_tsc_adjustment_strap,
       .fdtf_timestamp_valid,
       .fdtf_timestamp_value,
       .fdtf_force_ts,
       .ftrig_fabric_in,
       .atrig_fabric_in_ack,
       .atrig_fabric_out,
       .ftrig_fabric_out_ack,
       .dvp_paddr,
       .dvp_pprot,
       .dvp_psel,
       .dvp_penable,
       .dvp_pwrite,
       .dvp_pwdata,
       .dvp_pstrb,
       .dvp_pready,
       .dvp_pslverr,
       .dvp_prdata,
       .fdfx_powergood,
       .fdfx_earlyboot_debug_exit,
       .fdfx_policy_update,
       .fdfx_security_policy,
       .fdfx_debug_cap,
       .fdfx_debug_cap_valid);

   hqm_AW_clkbuf1 i_system_buf_hqm_clk_trunk
      (.a (prim_clk),
       .o (i_system_buf_hqm_clk_trunk_o));

   assign hqm_clk_enable                            = i_hqm_master_hqm_clk_enable;
   assign hqm_clk_rptr_rst_b                        = i_hqm_master_hqm_clk_rptr_rst_b;
   assign hqm_clk_trunk                             = i_system_buf_hqm_clk_trunk_o;
   assign hqm_clk_ungate                            = i_hqm_master_hqm_clk_ungate;
   assign hqm_gated_rst_b                           = hqm_gated_rst_b_mstr;
   assign hqm_proc_reset_done_sync_hqm              = i_hqm_master_hqm_proc_reset_done_sync_hqm;
   assign prim_clk_enable                           = i_hqm_sif_prim_clk_enable;
   assign prim_clk_ungate                           = i_hqm_sif_prim_clk_ungate;
   assign i_hqm_master_pgcb_isol_en_b               = pgcb_isol_en_b;


endmodule
