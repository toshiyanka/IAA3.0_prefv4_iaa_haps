### Tool : gds2def
### Version 14.1     Linux64
### Vendor : Apache Design, Inc. A Subsidiary of ANSYS, Inc. 
### Date : Jun 19 2014 02:20:56 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
MACRO c73p1rfshdxrom2048x32hb4img108_APACHECELL
 CLASS BLOCK ;
 ORIGIN 0 0 ;
 SIZE 75.432 BY 49.476 ;
 PIN iar[10]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 21.068 0.308 21.1 ;
 END
 END iar[10]
 PIN iar[0]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 21.754 0.308 21.786 ;
 END
 END iar[0]
 PIN iar[1]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 22.496 0.308 22.528 ;
 END
 END iar[1]
 PIN iar[2]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 23.126 0.308 23.158 ;
 END
 END iar[2]
 PIN iar[4]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 23.812 0.308 23.844 ;
 END
 END iar[4]
 PIN iar[3]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 24.442 0.308 24.474 ;
 END
 END iar[3]
 PIN iar[7]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 25.744 0.308 25.776 ;
 END
 END iar[7]
 PIN iar[6]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 26.43 0.308 26.462 ;
 END
 END iar[6]
 PIN iar[5]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 27.004 0.308 27.036 ;
 END
 END iar[5]
 PIN iar[9]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 27.802 0.308 27.834 ;
 END
 END iar[9]
 PIN iar[8]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 28.432 0.308 28.464 ;
 END
 END iar[8]
 PIN iren
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 25.184 0.308 25.216 ;
 END
 END iren
 PIN ickr
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 24.946 0.308 24.978 ;
 END
 END ickr
 PIN ipwreninb
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 48.718 0.308 48.75 ;
 END
 END ipwreninb
 PIN opwrenoutb
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 0.95 0.308 0.982 ;
 END
 END opwrenoutb
 PIN odout[0]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 1.062 0.308 1.094 ;
 END
 END odout[0]
 PIN odout[1]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 2.434 0.308 2.466 ;
 END
 END odout[1]
 PIN odout[2]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 3.694 0.308 3.726 ;
 END
 END odout[2]
 PIN odout[3]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 4.94 0.308 4.972 ;
 END
 END odout[3]
 PIN odout[4]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 6.088 0.308 6.12 ;
 END
 END odout[4]
 PIN odout[5]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 7.334 0.308 7.366 ;
 END
 END odout[5]
 PIN odout[6]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 8.594 0.308 8.626 ;
 END
 END odout[6]
 PIN odout[7]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 9.84 0.308 9.872 ;
 END
 END odout[7]
 PIN odout[8]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 11.212 0.308 11.244 ;
 END
 END odout[8]
 PIN odout[9]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 12.234 0.308 12.266 ;
 END
 END odout[9]
 PIN odout[10]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 13.494 0.308 13.526 ;
 END
 END odout[10]
 PIN odout[11]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 14.866 0.308 14.898 ;
 END
 END odout[11]
 PIN odout[12]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 16.224 0.308 16.256 ;
 END
 END odout[12]
 PIN odout[13]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 17.372 0.308 17.404 ;
 END
 END odout[13]
 PIN odout[14]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 18.618 0.308 18.65 ;
 END
 END odout[14]
 PIN odout[15]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 19.99 0.308 20.022 ;
 END
 END odout[15]
 PIN odout[16]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 29.342 0.308 29.374 ;
 END
 END odout[16]
 PIN odout[17]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 30.588 0.308 30.62 ;
 END
 END odout[17]
 PIN odout[18]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 31.624 0.308 31.656 ;
 END
 END odout[18]
 PIN odout[19]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 32.982 0.308 33.014 ;
 END
 END odout[19]
 PIN odout[20]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 34.354 0.308 34.386 ;
 END
 END odout[20]
 PIN odout[21]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 35.614 0.308 35.646 ;
 END
 END odout[21]
 PIN odout[22]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 36.748 0.308 36.78 ;
 END
 END odout[22]
 PIN odout[23]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 38.008 0.308 38.04 ;
 END
 END odout[23]
 PIN odout[24]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 39.254 0.308 39.286 ;
 END
 END odout[24]
 PIN odout[25]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 40.514 0.308 40.546 ;
 END
 END odout[25]
 PIN odout[26]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 41.76 0.308 41.792 ;
 END
 END odout[26]
 PIN odout[27]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 43.02 0.308 43.052 ;
 END
 END odout[27]
 PIN odout[28]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 44.154 0.308 44.186 ;
 END
 END odout[28]
 PIN odout[29]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 45.526 0.308 45.558 ;
 END
 END odout[29]
 PIN odout[30]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 46.898 0.308 46.93 ;
 END
 END odout[30]
 PIN odout[31]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER m4 ;
 RECT 0 48.144 0.308 48.176 ;
 END
 END odout[31]
 PIN vccd_1p0
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 2.978 0.43 3.178 ;
 END
 END vccd_1p0
 PIN vccd_1p0.gds1
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 1.013 1.542 1.213 ;
 END
 END vccd_1p0.gds1
 PIN vccd_1p0.gds2
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 1.022 5.202 1.222 ;
 END
 END vccd_1p0.gds2
 PIN vccd_1p0.gds3
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 2.273 1.542 2.473 ;
 END
 END vccd_1p0.gds3
 PIN vccd_1p0.gds4
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 4.793 1.542 4.993 ;
 END
 END vccd_1p0.gds4
 PIN vccd_1p0.gds5
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 4.6755 5.202 4.8755 ;
 END
 END vccd_1p0.gds5
 PIN vccd_1p0.gds6
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 3.089 0.548 3.289 ;
 END
 END vccd_1p0.gds6
 PIN vccd_1p0.gds7
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 3.0505 0.858 3.2505 ;
 END
 END vccd_1p0.gds7
 PIN vccd_1p0.gds8
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 2.888 1.362 3.088 ;
 END
 END vccd_1p0.gds8
 PIN vccd_1p0.gds9
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 3.106 1.782 3.306 ;
 END
 END vccd_1p0.gds9
 PIN vccd_1p0.gds10
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 2.987 1.218 3.187 ;
 END
 END vccd_1p0.gds10
 PIN vccd_1p0.gds11
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 3.533 1.542 3.733 ;
 END
 END vccd_1p0.gds11
 PIN vccd_1p0.gds12
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 3.4155 5.202 3.6155 ;
 END
 END vccd_1p0.gds12
 PIN vccd_1p0.gds13
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 3.061 1.962 3.261 ;
 END
 END vccd_1p0.gds13
 PIN vccd_1p0.gds14
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 2.9685 2.202 3.1685 ;
 END
 END vccd_1p0.gds14
 PIN vccd_1p0.gds15
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 3.0585 4.738 3.2585 ;
 END
 END vccd_1p0.gds15
 PIN vccd_1p0.gds16
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 3.0145 2.462 3.2145 ;
 END
 END vccd_1p0.gds16
 PIN vccd_1p0.gds17
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 3.007 2.622 3.207 ;
 END
 END vccd_1p0.gds17
 PIN vccd_1p0.gds18
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 3.007 1.09 3.207 ;
 END
 END vccd_1p0.gds18
 PIN vccd_1p0.gds19
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 2.8915 3.042 3.0915 ;
 END
 END vccd_1p0.gds19
 PIN vccd_1p0.gds20
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 3.02 2.882 3.22 ;
 END
 END vccd_1p0.gds20
 PIN vccd_1p0.gds21
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 2.98 3.39 3.18 ;
 END
 END vccd_1p0.gds21
 PIN vccd_1p0.gds22
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 3.016 3.262 3.216 ;
 END
 END vccd_1p0.gds22
 PIN vccd_1p0.gds23
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 2.1555 5.202 2.3555 ;
 END
 END vccd_1p0.gds23
 PIN vccd_1p0.gds24
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 3.059 3.666 3.259 ;
 END
 END vccd_1p0.gds24
 PIN vccd_1p0.gds25
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 3.0725 4.066 3.2725 ;
 END
 END vccd_1p0.gds25
 PIN vccd_1p0.gds26
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 3.0725 3.858 3.2725 ;
 END
 END vccd_1p0.gds26
 PIN vccd_1p0.gds27
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 3.02 4.258 3.22 ;
 END
 END vccd_1p0.gds27
 PIN vccd_1p0.gds28
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 3.058 4.546 3.258 ;
 END
 END vccd_1p0.gds28
 PIN vccd_1p0.gds29
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 3.082 5.01 3.282 ;
 END
 END vccd_1p0.gds29
 PIN vccd_1p0.gds30
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 4.34 1.228 4.396 1.428 ;
 RECT 4.76 1.204 4.816 1.404 ;
 RECT 5.096 1.228 5.152 1.428 ;
 RECT 4.34 2.488 4.396 2.688 ;
 RECT 4.76 2.464 4.816 2.664 ;
 RECT 5.096 2.488 5.152 2.688 ;
 RECT 4.34 3.748 4.396 3.948 ;
 RECT 4.76 3.724 4.816 3.924 ;
 RECT 5.096 3.748 5.152 3.948 ;
 RECT 4.34 5.008 4.396 5.208 ;
 RECT 4.76 4.984 4.816 5.184 ;
 RECT 5.096 5.008 5.152 5.208 ;
 RECT 3.584 4.8195 3.64 5.0195 ;
 RECT 4.172 4.9055 4.228 5.1055 ;
 RECT 4.928 4.862 4.984 5.062 ;
 RECT 3.584 3.5595 3.64 3.7595 ;
 RECT 4.172 3.6455 4.228 3.8455 ;
 RECT 4.928 3.602 4.984 3.802 ;
 RECT 3.584 2.2995 3.64 2.4995 ;
 RECT 4.172 2.3855 4.228 2.5855 ;
 RECT 4.928 2.342 4.984 2.542 ;
 RECT 3.584 1.0395 3.64 1.2395 ;
 RECT 4.172 1.1255 4.228 1.3255 ;
 RECT 4.928 1.082 4.984 1.282 ;
 END
 END vccd_1p0.gds30
 PIN vccd_1p0.gds31
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 3.0725 6.838 3.2725 ;
 END
 END vccd_1p0.gds31
 PIN vccd_1p0.gds32
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 3.082 6.05 3.282 ;
 END
 END vccd_1p0.gds32
 PIN vccd_1p0.gds33
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.754 3.02 5.794 3.22 ;
 END
 END vccd_1p0.gds33
 PIN vccd_1p0.gds34
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 3.109 6.306 3.309 ;
 END
 END vccd_1p0.gds34
 PIN vccd_1p0.gds35
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 3.0725 5.41 3.2725 ;
 END
 END vccd_1p0.gds35
 PIN vccd_1p0.gds36
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 3.0725 5.922 3.2725 ;
 END
 END vccd_1p0.gds36
 PIN vccd_1p0.gds37
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 2.962 5.602 3.162 ;
 END
 END vccd_1p0.gds37
 PIN vccd_1p0.gds38
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 2.999 6.582 3.199 ;
 END
 END vccd_1p0.gds38
 PIN vccd_1p0.gds39
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.6 4.9055 5.656 5.1055 ;
 RECT 5.264 4.9055 5.32 5.1055 ;
 RECT 5.432 4.8195 5.488 5.0195 ;
 RECT 5.936 4.8195 5.992 5.0195 ;
 RECT 5.768 4.8195 5.824 5.0195 ;
 RECT 6.44 4.834 6.496 5.034 ;
 RECT 6.272 4.8195 6.328 5.0195 ;
 RECT 6.104 5.008 6.16 5.208 ;
 RECT 5.6 3.6455 5.656 3.8455 ;
 RECT 5.264 3.6455 5.32 3.8455 ;
 RECT 5.432 3.5595 5.488 3.7595 ;
 RECT 5.936 3.5595 5.992 3.7595 ;
 RECT 5.768 3.5595 5.824 3.7595 ;
 RECT 6.44 3.574 6.496 3.774 ;
 RECT 6.272 3.5595 6.328 3.7595 ;
 RECT 6.104 3.748 6.16 3.948 ;
 RECT 5.6 2.3855 5.656 2.5855 ;
 RECT 5.264 2.3855 5.32 2.5855 ;
 RECT 5.432 2.2995 5.488 2.4995 ;
 RECT 5.936 2.2995 5.992 2.4995 ;
 RECT 5.768 2.2995 5.824 2.4995 ;
 RECT 6.44 2.314 6.496 2.514 ;
 RECT 6.272 2.2995 6.328 2.4995 ;
 RECT 6.104 2.488 6.16 2.688 ;
 RECT 5.6 1.1255 5.656 1.3255 ;
 RECT 5.264 1.1255 5.32 1.3255 ;
 RECT 5.432 1.0395 5.488 1.2395 ;
 RECT 5.936 1.0395 5.992 1.2395 ;
 RECT 5.768 1.0395 5.824 1.2395 ;
 RECT 6.44 1.054 6.496 1.254 ;
 RECT 6.272 1.0395 6.328 1.2395 ;
 RECT 6.104 1.228 6.16 1.428 ;
 END
 END vccd_1p0.gds39
 PIN vccd_1p0.gds40
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 1.36 13.978 1.56 ;
 END
 END vccd_1p0.gds40
 PIN vccd_1p0.gds41
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 2.62 13.978 2.82 ;
 END
 END vccd_1p0.gds41
 PIN vccd_1p0.gds42
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 3.88 13.978 4.08 ;
 END
 END vccd_1p0.gds42
 PIN vccd_1p0.gds43
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 5.14 14.398 5.34 ;
 END
 END vccd_1p0.gds43
 PIN vccd_1p0.gds44
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 5.2675 14.934 5.4675 ;
 END
 END vccd_1p0.gds44
 PIN vccd_1p0.gds45
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 3.88 14.398 4.08 ;
 END
 END vccd_1p0.gds45
 PIN vccd_1p0.gds46
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 4.0075 14.934 4.2075 ;
 END
 END vccd_1p0.gds46
 PIN vccd_1p0.gds47
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 2.62 14.398 2.82 ;
 END
 END vccd_1p0.gds47
 PIN vccd_1p0.gds48
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 2.7475 14.934 2.9475 ;
 END
 END vccd_1p0.gds48
 PIN vccd_1p0.gds49
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 1.36 14.398 1.56 ;
 END
 END vccd_1p0.gds49
 PIN vccd_1p0.gds50
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 1.4875 14.934 1.6875 ;
 END
 END vccd_1p0.gds50
 PIN vccd_1p0.gds51
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 3.072 14.742 3.272 ;
 END
 END vccd_1p0.gds51
 PIN vccd_1p0.gds52
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 5.14 13.978 5.34 ;
 END
 END vccd_1p0.gds52
 PIN vccd_1p0.gds53
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 2.82 13.738 3.02 ;
 END
 END vccd_1p0.gds53
 PIN vccd_1p0.gds54
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 3.02 12.898 3.22 ;
 END
 END vccd_1p0.gds54
 PIN vccd_1p0.gds55
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 2.8975 13.138 3.0975 ;
 END
 END vccd_1p0.gds55
 PIN vccd_1p0.gds56
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 3.016 12.654 3.216 ;
 END
 END vccd_1p0.gds56
 PIN vccd_1p0.gds57
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 2.9745 12.526 3.1745 ;
 END
 END vccd_1p0.gds57
 PIN vccd_1p0.gds58
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 1.424 16.226 1.624 ;
 END
 END vccd_1p0.gds58
 PIN vccd_1p0.gds59
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 5.204 16.226 5.404 ;
 END
 END vccd_1p0.gds59
 PIN vccd_1p0.gds60
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 3.944 16.226 4.144 ;
 END
 END vccd_1p0.gds60
 PIN vccd_1p0.gds61
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 2.684 16.226 2.884 ;
 END
 END vccd_1p0.gds61
 PIN vccd_1p0.gds62
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 3.054 15.742 3.254 ;
 END
 END vccd_1p0.gds62
 PIN vccd_1p0.gds63
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 3.072 15.29 3.272 ;
 END
 END vccd_1p0.gds63
 PIN vccd_1p0.gds64
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 2.9985 17.574 3.1985 ;
 END
 END vccd_1p0.gds64
 PIN vccd_1p0.gds65
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 2.9235 17.154 3.1235 ;
 END
 END vccd_1p0.gds65
 PIN vccd_1p0.gds66
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 3.02 17.734 3.22 ;
 END
 END vccd_1p0.gds66
 PIN vccd_1p0.gds67
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 3.054 15.498 3.254 ;
 END
 END vccd_1p0.gds67
 PIN vccd_1p0.gds68
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 3.016 17.962 3.216 ;
 END
 END vccd_1p0.gds68
 PIN vccd_1p0.gds69
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 2.9745 18.09 3.1745 ;
 END
 END vccd_1p0.gds69
 PIN vccd_1p0.gds70
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 2.9785 23.842 3.1785 ;
 END
 END vccd_1p0.gds70
 PIN vccd_1p0.gds71
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 3.02 29.95 3.22 ;
 END
 END vccd_1p0.gds71
 PIN vccd_1p0.gds72
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 3.016 29.706 3.216 ;
 END
 END vccd_1p0.gds72
 PIN vccd_1p0.gds73
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 2.9745 29.578 3.1745 ;
 END
 END vccd_1p0.gds73
 PIN vccd_1p0.gds74
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 1.424 33.278 1.624 ;
 END
 END vccd_1p0.gds74
 PIN vccd_1p0.gds75
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 1.36 31.45 1.56 ;
 END
 END vccd_1p0.gds75
 PIN vccd_1p0.gds76
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 2.684 33.278 2.884 ;
 END
 END vccd_1p0.gds76
 PIN vccd_1p0.gds77
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 2.62 31.45 2.82 ;
 END
 END vccd_1p0.gds77
 PIN vccd_1p0.gds78
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 3.944 33.278 4.144 ;
 END
 END vccd_1p0.gds78
 PIN vccd_1p0.gds79
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 1.36 31.03 1.56 ;
 END
 END vccd_1p0.gds79
 PIN vccd_1p0.gds80
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 2.62 31.03 2.82 ;
 END
 END vccd_1p0.gds80
 PIN vccd_1p0.gds81
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 5.14 31.03 5.34 ;
 END
 END vccd_1p0.gds81
 PIN vccd_1p0.gds82
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 3.88 31.03 4.08 ;
 END
 END vccd_1p0.gds82
 PIN vccd_1p0.gds83
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 2.82 30.79 3.02 ;
 END
 END vccd_1p0.gds83
 PIN vccd_1p0.gds84
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 2.8975 30.19 3.0975 ;
 END
 END vccd_1p0.gds84
 PIN vccd_1p0.gds85
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 5.204 33.278 5.404 ;
 END
 END vccd_1p0.gds85
 PIN vccd_1p0.gds86
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 5.14 31.45 5.34 ;
 END
 END vccd_1p0.gds86
 PIN vccd_1p0.gds87
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 5.2675 31.986 5.4675 ;
 END
 END vccd_1p0.gds87
 PIN vccd_1p0.gds88
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 3.072 32.342 3.272 ;
 END
 END vccd_1p0.gds88
 PIN vccd_1p0.gds89
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 3.072 31.794 3.272 ;
 END
 END vccd_1p0.gds89
 PIN vccd_1p0.gds90
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 3.88 31.45 4.08 ;
 END
 END vccd_1p0.gds90
 PIN vccd_1p0.gds91
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 4.0075 31.986 4.2075 ;
 END
 END vccd_1p0.gds91
 PIN vccd_1p0.gds92
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 2.9985 34.626 3.1985 ;
 END
 END vccd_1p0.gds92
 PIN vccd_1p0.gds93
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 2.9745 35.142 3.1745 ;
 END
 END vccd_1p0.gds93
 PIN vccd_1p0.gds94
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 3.016 35.014 3.216 ;
 END
 END vccd_1p0.gds94
 PIN vccd_1p0.gds95
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 2.9235 34.206 3.1235 ;
 END
 END vccd_1p0.gds95
 PIN vccd_1p0.gds96
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 2.7475 31.986 2.9475 ;
 END
 END vccd_1p0.gds96
 PIN vccd_1p0.gds97
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 3.054 32.794 3.254 ;
 END
 END vccd_1p0.gds97
 PIN vccd_1p0.gds98
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 3.054 32.55 3.254 ;
 END
 END vccd_1p0.gds98
 PIN vccd_1p0.gds99
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 1.4875 31.986 1.6875 ;
 END
 END vccd_1p0.gds99
 PIN vccd_1p0.gds100
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 3.02 34.786 3.22 ;
 END
 END vccd_1p0.gds100
 PIN vccd_1p0.gds101
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 2.9785 40.894 3.1785 ;
 END
 END vccd_1p0.gds101
 PIN vccd_1p0.gds102
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 1.36 48.082 1.56 ;
 END
 END vccd_1p0.gds102
 PIN vccd_1p0.gds103
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 2.62 48.082 2.82 ;
 END
 END vccd_1p0.gds103
 PIN vccd_1p0.gds104
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 3.88 48.082 4.08 ;
 END
 END vccd_1p0.gds104
 PIN vccd_1p0.gds105
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 5.14 48.082 5.34 ;
 END
 END vccd_1p0.gds105
 PIN vccd_1p0.gds106
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 1.36 48.502 1.56 ;
 END
 END vccd_1p0.gds106
 PIN vccd_1p0.gds107
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 2.62 48.502 2.82 ;
 END
 END vccd_1p0.gds107
 PIN vccd_1p0.gds108
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 2.82 47.842 3.02 ;
 END
 END vccd_1p0.gds108
 PIN vccd_1p0.gds109
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 2.8975 47.242 3.0975 ;
 END
 END vccd_1p0.gds109
 PIN vccd_1p0.gds110
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 5.14 48.502 5.34 ;
 END
 END vccd_1p0.gds110
 PIN vccd_1p0.gds111
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 5.2675 49.038 5.4675 ;
 END
 END vccd_1p0.gds111
 PIN vccd_1p0.gds112
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 3.072 49.394 3.272 ;
 END
 END vccd_1p0.gds112
 PIN vccd_1p0.gds113
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 3.072 48.846 3.272 ;
 END
 END vccd_1p0.gds113
 PIN vccd_1p0.gds114
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 3.88 48.502 4.08 ;
 END
 END vccd_1p0.gds114
 PIN vccd_1p0.gds115
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 4.0075 49.038 4.2075 ;
 END
 END vccd_1p0.gds115
 PIN vccd_1p0.gds116
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 2.7475 49.038 2.9475 ;
 END
 END vccd_1p0.gds116
 PIN vccd_1p0.gds117
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 3.054 49.846 3.254 ;
 END
 END vccd_1p0.gds117
 PIN vccd_1p0.gds118
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 3.054 49.602 3.254 ;
 END
 END vccd_1p0.gds118
 PIN vccd_1p0.gds119
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 1.4875 49.038 1.6875 ;
 END
 END vccd_1p0.gds119
 PIN vccd_1p0.gds120
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 3.02 47.002 3.22 ;
 END
 END vccd_1p0.gds120
 PIN vccd_1p0.gds121
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 3.016 46.758 3.216 ;
 END
 END vccd_1p0.gds121
 PIN vccd_1p0.gds122
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 2.9745 46.63 3.1745 ;
 END
 END vccd_1p0.gds122
 PIN vccd_1p0.gds123
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 1.424 50.33 1.624 ;
 END
 END vccd_1p0.gds123
 PIN vccd_1p0.gds124
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 2.684 50.33 2.884 ;
 END
 END vccd_1p0.gds124
 PIN vccd_1p0.gds125
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 3.944 50.33 4.144 ;
 END
 END vccd_1p0.gds125
 PIN vccd_1p0.gds126
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 5.204 50.33 5.404 ;
 END
 END vccd_1p0.gds126
 PIN vccd_1p0.gds127
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 2.9985 51.678 3.1985 ;
 END
 END vccd_1p0.gds127
 PIN vccd_1p0.gds128
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 2.9745 52.194 3.1745 ;
 END
 END vccd_1p0.gds128
 PIN vccd_1p0.gds129
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 3.016 52.066 3.216 ;
 END
 END vccd_1p0.gds129
 PIN vccd_1p0.gds130
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 2.9235 51.258 3.1235 ;
 END
 END vccd_1p0.gds130
 PIN vccd_1p0.gds131
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 3.02 51.838 3.22 ;
 END
 END vccd_1p0.gds131
 PIN vccd_1p0.gds132
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 2.9785 57.946 3.1785 ;
 END
 END vccd_1p0.gds132
 PIN vccd_1p0.gds133
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 1.36 65.134 1.56 ;
 END
 END vccd_1p0.gds133
 PIN vccd_1p0.gds134
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 2.62 65.134 2.82 ;
 END
 END vccd_1p0.gds134
 PIN vccd_1p0.gds135
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 3.88 65.134 4.08 ;
 END
 END vccd_1p0.gds135
 PIN vccd_1p0.gds136
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 5.14 65.134 5.34 ;
 END
 END vccd_1p0.gds136
 PIN vccd_1p0.gds137
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 2.82 64.894 3.02 ;
 END
 END vccd_1p0.gds137
 PIN vccd_1p0.gds138
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 2.8975 64.294 3.0975 ;
 END
 END vccd_1p0.gds138
 PIN vccd_1p0.gds139
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 3.02 64.054 3.22 ;
 END
 END vccd_1p0.gds139
 PIN vccd_1p0.gds140
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 3.016 63.81 3.216 ;
 END
 END vccd_1p0.gds140
 PIN vccd_1p0.gds141
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 2.9745 63.682 3.1745 ;
 END
 END vccd_1p0.gds141
 PIN vccd_1p0.gds142
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 1.424 67.382 1.624 ;
 END
 END vccd_1p0.gds142
 PIN vccd_1p0.gds143
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 1.36 65.554 1.56 ;
 END
 END vccd_1p0.gds143
 PIN vccd_1p0.gds144
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 2.684 67.382 2.884 ;
 END
 END vccd_1p0.gds144
 PIN vccd_1p0.gds145
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 2.62 65.554 2.82 ;
 END
 END vccd_1p0.gds145
 PIN vccd_1p0.gds146
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 3.944 67.382 4.144 ;
 END
 END vccd_1p0.gds146
 PIN vccd_1p0.gds147
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 5.204 67.382 5.404 ;
 END
 END vccd_1p0.gds147
 PIN vccd_1p0.gds148
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 5.14 65.554 5.34 ;
 END
 END vccd_1p0.gds148
 PIN vccd_1p0.gds149
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 5.2675 66.09 5.4675 ;
 END
 END vccd_1p0.gds149
 PIN vccd_1p0.gds150
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 3.072 66.446 3.272 ;
 END
 END vccd_1p0.gds150
 PIN vccd_1p0.gds151
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 3.072 65.898 3.272 ;
 END
 END vccd_1p0.gds151
 PIN vccd_1p0.gds152
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 3.88 65.554 4.08 ;
 END
 END vccd_1p0.gds152
 PIN vccd_1p0.gds153
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 4.0075 66.09 4.2075 ;
 END
 END vccd_1p0.gds153
 PIN vccd_1p0.gds154
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 2.9985 68.73 3.1985 ;
 END
 END vccd_1p0.gds154
 PIN vccd_1p0.gds155
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 2.9745 69.246 3.1745 ;
 END
 END vccd_1p0.gds155
 PIN vccd_1p0.gds156
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 3.016 69.118 3.216 ;
 END
 END vccd_1p0.gds156
 PIN vccd_1p0.gds157
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 2.9235 68.31 3.1235 ;
 END
 END vccd_1p0.gds157
 PIN vccd_1p0.gds158
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 2.7475 66.09 2.9475 ;
 END
 END vccd_1p0.gds158
 PIN vccd_1p0.gds159
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 3.054 66.898 3.254 ;
 END
 END vccd_1p0.gds159
 PIN vccd_1p0.gds160
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 3.054 66.654 3.254 ;
 END
 END vccd_1p0.gds160
 PIN vccd_1p0.gds161
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 1.4875 66.09 1.6875 ;
 END
 END vccd_1p0.gds161
 PIN vccd_1p0.gds162
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 3.02 68.89 3.22 ;
 END
 END vccd_1p0.gds162
 PIN vccd_1p0.gds163
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 8.018 0.43 8.218 ;
 END
 END vccd_1p0.gds163
 PIN vccd_1p0.gds164
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 9.833 1.542 10.033 ;
 END
 END vccd_1p0.gds164
 PIN vccd_1p0.gds165
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 9.7155 5.202 9.9155 ;
 END
 END vccd_1p0.gds165
 PIN vccd_1p0.gds166
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 8.573 1.542 8.773 ;
 END
 END vccd_1p0.gds166
 PIN vccd_1p0.gds167
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 8.4555 5.202 8.6555 ;
 END
 END vccd_1p0.gds167
 PIN vccd_1p0.gds168
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 7.313 1.542 7.513 ;
 END
 END vccd_1p0.gds168
 PIN vccd_1p0.gds169
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 7.1955 5.202 7.3955 ;
 END
 END vccd_1p0.gds169
 PIN vccd_1p0.gds170
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 6.053 1.542 6.253 ;
 END
 END vccd_1p0.gds170
 PIN vccd_1p0.gds171
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 5.9355 5.202 6.1355 ;
 END
 END vccd_1p0.gds171
 PIN vccd_1p0.gds172
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 8.129 0.548 8.329 ;
 END
 END vccd_1p0.gds172
 PIN vccd_1p0.gds173
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 8.0905 0.858 8.2905 ;
 END
 END vccd_1p0.gds173
 PIN vccd_1p0.gds174
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 7.928 1.362 8.128 ;
 END
 END vccd_1p0.gds174
 PIN vccd_1p0.gds175
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 8.146 1.782 8.346 ;
 END
 END vccd_1p0.gds175
 PIN vccd_1p0.gds176
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 8.027 1.218 8.227 ;
 END
 END vccd_1p0.gds176
 PIN vccd_1p0.gds177
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 8.101 1.962 8.301 ;
 END
 END vccd_1p0.gds177
 PIN vccd_1p0.gds178
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 8.0085 2.202 8.2085 ;
 END
 END vccd_1p0.gds178
 PIN vccd_1p0.gds179
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 8.0985 4.738 8.2985 ;
 END
 END vccd_1p0.gds179
 PIN vccd_1p0.gds180
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 8.0545 2.462 8.2545 ;
 END
 END vccd_1p0.gds180
 PIN vccd_1p0.gds181
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 8.047 2.622 8.247 ;
 END
 END vccd_1p0.gds181
 PIN vccd_1p0.gds182
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 8.047 1.09 8.247 ;
 END
 END vccd_1p0.gds182
 PIN vccd_1p0.gds183
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 7.9315 3.042 8.1315 ;
 END
 END vccd_1p0.gds183
 PIN vccd_1p0.gds184
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 8.06 2.882 8.26 ;
 END
 END vccd_1p0.gds184
 PIN vccd_1p0.gds185
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 8.02 3.39 8.22 ;
 END
 END vccd_1p0.gds185
 PIN vccd_1p0.gds186
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 8.056 3.262 8.256 ;
 END
 END vccd_1p0.gds186
 PIN vccd_1p0.gds187
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 8.099 3.666 8.299 ;
 END
 END vccd_1p0.gds187
 PIN vccd_1p0.gds188
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 8.1125 4.066 8.3125 ;
 END
 END vccd_1p0.gds188
 PIN vccd_1p0.gds189
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 8.1125 3.858 8.3125 ;
 END
 END vccd_1p0.gds189
 PIN vccd_1p0.gds190
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 8.06 4.258 8.26 ;
 END
 END vccd_1p0.gds190
 PIN vccd_1p0.gds191
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 8.098 4.546 8.298 ;
 END
 END vccd_1p0.gds191
 PIN vccd_1p0.gds192
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 8.122 5.01 8.322 ;
 END
 END vccd_1p0.gds192
 PIN vccd_1p0.gds193
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 4.34 6.268 4.396 6.468 ;
 RECT 4.76 6.244 4.816 6.444 ;
 RECT 5.096 6.268 5.152 6.468 ;
 RECT 4.34 7.528 4.396 7.728 ;
 RECT 4.76 7.504 4.816 7.704 ;
 RECT 5.096 7.528 5.152 7.728 ;
 RECT 4.34 8.788 4.396 8.988 ;
 RECT 4.76 8.764 4.816 8.964 ;
 RECT 5.096 8.788 5.152 8.988 ;
 RECT 4.34 10.048 4.396 10.248 ;
 RECT 4.76 10.024 4.816 10.224 ;
 RECT 5.096 10.048 5.152 10.248 ;
 RECT 3.584 9.8595 3.64 10.0595 ;
 RECT 4.172 9.9455 4.228 10.1455 ;
 RECT 4.928 9.902 4.984 10.102 ;
 RECT 3.584 8.5995 3.64 8.7995 ;
 RECT 4.172 8.6855 4.228 8.8855 ;
 RECT 4.928 8.642 4.984 8.842 ;
 RECT 3.584 7.3395 3.64 7.5395 ;
 RECT 4.172 7.4255 4.228 7.6255 ;
 RECT 4.928 7.382 4.984 7.582 ;
 RECT 3.584 6.0795 3.64 6.2795 ;
 RECT 4.172 6.1655 4.228 6.3655 ;
 RECT 4.928 6.122 4.984 6.322 ;
 END
 END vccd_1p0.gds193
 PIN vccd_1p0.gds194
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 8.1125 6.838 8.3125 ;
 END
 END vccd_1p0.gds194
 PIN vccd_1p0.gds195
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 8.122 6.05 8.322 ;
 END
 END vccd_1p0.gds195
 PIN vccd_1p0.gds196
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.754 8.06 5.794 8.26 ;
 END
 END vccd_1p0.gds196
 PIN vccd_1p0.gds197
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 8.149 6.306 8.349 ;
 END
 END vccd_1p0.gds197
 PIN vccd_1p0.gds198
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 8.1125 5.41 8.3125 ;
 END
 END vccd_1p0.gds198
 PIN vccd_1p0.gds199
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 8.1125 5.922 8.3125 ;
 END
 END vccd_1p0.gds199
 PIN vccd_1p0.gds200
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 8.002 5.602 8.202 ;
 END
 END vccd_1p0.gds200
 PIN vccd_1p0.gds201
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 8.039 6.582 8.239 ;
 END
 END vccd_1p0.gds201
 PIN vccd_1p0.gds202
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.6 9.9455 5.656 10.1455 ;
 RECT 5.264 9.9455 5.32 10.1455 ;
 RECT 5.432 9.8595 5.488 10.0595 ;
 RECT 5.936 9.8595 5.992 10.0595 ;
 RECT 5.768 9.8595 5.824 10.0595 ;
 RECT 6.44 9.874 6.496 10.074 ;
 RECT 6.272 9.8595 6.328 10.0595 ;
 RECT 6.104 10.048 6.16 10.248 ;
 RECT 5.6 8.6855 5.656 8.8855 ;
 RECT 5.264 8.6855 5.32 8.8855 ;
 RECT 5.432 8.5995 5.488 8.7995 ;
 RECT 5.936 8.5995 5.992 8.7995 ;
 RECT 5.768 8.5995 5.824 8.7995 ;
 RECT 6.44 8.614 6.496 8.814 ;
 RECT 6.272 8.5995 6.328 8.7995 ;
 RECT 6.104 8.788 6.16 8.988 ;
 RECT 5.6 7.4255 5.656 7.6255 ;
 RECT 5.264 7.4255 5.32 7.6255 ;
 RECT 5.432 7.3395 5.488 7.5395 ;
 RECT 5.936 7.3395 5.992 7.5395 ;
 RECT 5.768 7.3395 5.824 7.5395 ;
 RECT 6.44 7.354 6.496 7.554 ;
 RECT 6.272 7.3395 6.328 7.5395 ;
 RECT 6.104 7.528 6.16 7.728 ;
 RECT 5.6 6.1655 5.656 6.3655 ;
 RECT 5.264 6.1655 5.32 6.3655 ;
 RECT 5.432 6.0795 5.488 6.2795 ;
 RECT 5.936 6.0795 5.992 6.2795 ;
 RECT 5.768 6.0795 5.824 6.2795 ;
 RECT 6.44 6.094 6.496 6.294 ;
 RECT 6.272 6.0795 6.328 6.2795 ;
 RECT 6.104 6.268 6.16 6.468 ;
 END
 END vccd_1p0.gds202
 PIN vccd_1p0.gds203
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 6.4 13.978 6.6 ;
 END
 END vccd_1p0.gds203
 PIN vccd_1p0.gds204
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 7.66 13.978 7.86 ;
 END
 END vccd_1p0.gds204
 PIN vccd_1p0.gds205
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 8.92 13.978 9.12 ;
 END
 END vccd_1p0.gds205
 PIN vccd_1p0.gds206
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 10.18 13.978 10.38 ;
 END
 END vccd_1p0.gds206
 PIN vccd_1p0.gds207
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 10.18 14.398 10.38 ;
 END
 END vccd_1p0.gds207
 PIN vccd_1p0.gds208
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 10.3075 14.934 10.5075 ;
 END
 END vccd_1p0.gds208
 PIN vccd_1p0.gds209
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 8.92 14.398 9.12 ;
 END
 END vccd_1p0.gds209
 PIN vccd_1p0.gds210
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 9.0475 14.934 9.2475 ;
 END
 END vccd_1p0.gds210
 PIN vccd_1p0.gds211
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 7.66 14.398 7.86 ;
 END
 END vccd_1p0.gds211
 PIN vccd_1p0.gds212
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 7.7875 14.934 7.9875 ;
 END
 END vccd_1p0.gds212
 PIN vccd_1p0.gds213
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 6.4 14.398 6.6 ;
 END
 END vccd_1p0.gds213
 PIN vccd_1p0.gds214
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 6.5275 14.934 6.7275 ;
 END
 END vccd_1p0.gds214
 PIN vccd_1p0.gds215
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 8.112 14.742 8.312 ;
 END
 END vccd_1p0.gds215
 PIN vccd_1p0.gds216
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 7.86 13.738 8.06 ;
 END
 END vccd_1p0.gds216
 PIN vccd_1p0.gds217
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 8.06 12.898 8.26 ;
 END
 END vccd_1p0.gds217
 PIN vccd_1p0.gds218
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 7.9375 13.138 8.1375 ;
 END
 END vccd_1p0.gds218
 PIN vccd_1p0.gds219
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 8.056 12.654 8.256 ;
 END
 END vccd_1p0.gds219
 PIN vccd_1p0.gds220
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 8.0145 12.526 8.2145 ;
 END
 END vccd_1p0.gds220
 PIN vccd_1p0.gds221
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 10.244 16.226 10.444 ;
 END
 END vccd_1p0.gds221
 PIN vccd_1p0.gds222
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 8.984 16.226 9.184 ;
 END
 END vccd_1p0.gds222
 PIN vccd_1p0.gds223
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 7.724 16.226 7.924 ;
 END
 END vccd_1p0.gds223
 PIN vccd_1p0.gds224
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 6.464 16.226 6.664 ;
 END
 END vccd_1p0.gds224
 PIN vccd_1p0.gds225
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 8.094 15.742 8.294 ;
 END
 END vccd_1p0.gds225
 PIN vccd_1p0.gds226
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 8.112 15.29 8.312 ;
 END
 END vccd_1p0.gds226
 PIN vccd_1p0.gds227
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 8.0385 17.574 8.2385 ;
 END
 END vccd_1p0.gds227
 PIN vccd_1p0.gds228
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 7.9635 17.154 8.1635 ;
 END
 END vccd_1p0.gds228
 PIN vccd_1p0.gds229
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 8.06 17.734 8.26 ;
 END
 END vccd_1p0.gds229
 PIN vccd_1p0.gds230
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 8.094 15.498 8.294 ;
 END
 END vccd_1p0.gds230
 PIN vccd_1p0.gds231
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 8.056 17.962 8.256 ;
 END
 END vccd_1p0.gds231
 PIN vccd_1p0.gds232
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 8.0145 18.09 8.2145 ;
 END
 END vccd_1p0.gds232
 PIN vccd_1p0.gds233
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 8.0185 23.842 8.2185 ;
 END
 END vccd_1p0.gds233
 PIN vccd_1p0.gds234
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 8.06 29.95 8.26 ;
 END
 END vccd_1p0.gds234
 PIN vccd_1p0.gds235
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 8.056 29.706 8.256 ;
 END
 END vccd_1p0.gds235
 PIN vccd_1p0.gds236
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 8.0145 29.578 8.2145 ;
 END
 END vccd_1p0.gds236
 PIN vccd_1p0.gds237
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 10.18 31.03 10.38 ;
 END
 END vccd_1p0.gds237
 PIN vccd_1p0.gds238
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 8.92 31.03 9.12 ;
 END
 END vccd_1p0.gds238
 PIN vccd_1p0.gds239
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 6.464 33.278 6.664 ;
 END
 END vccd_1p0.gds239
 PIN vccd_1p0.gds240
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 6.4 31.45 6.6 ;
 END
 END vccd_1p0.gds240
 PIN vccd_1p0.gds241
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 6.5275 31.986 6.7275 ;
 END
 END vccd_1p0.gds241
 PIN vccd_1p0.gds242
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 7.724 33.278 7.924 ;
 END
 END vccd_1p0.gds242
 PIN vccd_1p0.gds243
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 7.66 31.45 7.86 ;
 END
 END vccd_1p0.gds243
 PIN vccd_1p0.gds244
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 7.7875 31.986 7.9875 ;
 END
 END vccd_1p0.gds244
 PIN vccd_1p0.gds245
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 8.984 33.278 9.184 ;
 END
 END vccd_1p0.gds245
 PIN vccd_1p0.gds246
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 8.92 31.45 9.12 ;
 END
 END vccd_1p0.gds246
 PIN vccd_1p0.gds247
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 9.0475 31.986 9.2475 ;
 END
 END vccd_1p0.gds247
 PIN vccd_1p0.gds248
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 10.244 33.278 10.444 ;
 END
 END vccd_1p0.gds248
 PIN vccd_1p0.gds249
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 10.18 31.45 10.38 ;
 END
 END vccd_1p0.gds249
 PIN vccd_1p0.gds250
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 10.3075 31.986 10.5075 ;
 END
 END vccd_1p0.gds250
 PIN vccd_1p0.gds251
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 7.66 31.03 7.86 ;
 END
 END vccd_1p0.gds251
 PIN vccd_1p0.gds252
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 6.4 31.03 6.6 ;
 END
 END vccd_1p0.gds252
 PIN vccd_1p0.gds253
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 7.86 30.79 8.06 ;
 END
 END vccd_1p0.gds253
 PIN vccd_1p0.gds254
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 7.9375 30.19 8.1375 ;
 END
 END vccd_1p0.gds254
 PIN vccd_1p0.gds255
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 8.112 32.342 8.312 ;
 END
 END vccd_1p0.gds255
 PIN vccd_1p0.gds256
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 8.112 31.794 8.312 ;
 END
 END vccd_1p0.gds256
 PIN vccd_1p0.gds257
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 8.0385 34.626 8.2385 ;
 END
 END vccd_1p0.gds257
 PIN vccd_1p0.gds258
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 8.0145 35.142 8.2145 ;
 END
 END vccd_1p0.gds258
 PIN vccd_1p0.gds259
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 8.056 35.014 8.256 ;
 END
 END vccd_1p0.gds259
 PIN vccd_1p0.gds260
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 7.9635 34.206 8.1635 ;
 END
 END vccd_1p0.gds260
 PIN vccd_1p0.gds261
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 8.094 32.794 8.294 ;
 END
 END vccd_1p0.gds261
 PIN vccd_1p0.gds262
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 8.094 32.55 8.294 ;
 END
 END vccd_1p0.gds262
 PIN vccd_1p0.gds263
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 8.06 34.786 8.26 ;
 END
 END vccd_1p0.gds263
 PIN vccd_1p0.gds264
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 8.0185 40.894 8.2185 ;
 END
 END vccd_1p0.gds264
 PIN vccd_1p0.gds265
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 6.4 48.082 6.6 ;
 END
 END vccd_1p0.gds265
 PIN vccd_1p0.gds266
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 7.66 48.082 7.86 ;
 END
 END vccd_1p0.gds266
 PIN vccd_1p0.gds267
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 8.92 48.082 9.12 ;
 END
 END vccd_1p0.gds267
 PIN vccd_1p0.gds268
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 10.18 48.082 10.38 ;
 END
 END vccd_1p0.gds268
 PIN vccd_1p0.gds269
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 10.18 48.502 10.38 ;
 END
 END vccd_1p0.gds269
 PIN vccd_1p0.gds270
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 10.3075 49.038 10.5075 ;
 END
 END vccd_1p0.gds270
 PIN vccd_1p0.gds271
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 8.92 48.502 9.12 ;
 END
 END vccd_1p0.gds271
 PIN vccd_1p0.gds272
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 9.0475 49.038 9.2475 ;
 END
 END vccd_1p0.gds272
 PIN vccd_1p0.gds273
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 7.66 48.502 7.86 ;
 END
 END vccd_1p0.gds273
 PIN vccd_1p0.gds274
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 7.7875 49.038 7.9875 ;
 END
 END vccd_1p0.gds274
 PIN vccd_1p0.gds275
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 6.4 48.502 6.6 ;
 END
 END vccd_1p0.gds275
 PIN vccd_1p0.gds276
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 6.5275 49.038 6.7275 ;
 END
 END vccd_1p0.gds276
 PIN vccd_1p0.gds277
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 7.86 47.842 8.06 ;
 END
 END vccd_1p0.gds277
 PIN vccd_1p0.gds278
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 7.9375 47.242 8.1375 ;
 END
 END vccd_1p0.gds278
 PIN vccd_1p0.gds279
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 8.112 49.394 8.312 ;
 END
 END vccd_1p0.gds279
 PIN vccd_1p0.gds280
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 8.112 48.846 8.312 ;
 END
 END vccd_1p0.gds280
 PIN vccd_1p0.gds281
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 8.094 49.846 8.294 ;
 END
 END vccd_1p0.gds281
 PIN vccd_1p0.gds282
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 8.094 49.602 8.294 ;
 END
 END vccd_1p0.gds282
 PIN vccd_1p0.gds283
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 8.06 47.002 8.26 ;
 END
 END vccd_1p0.gds283
 PIN vccd_1p0.gds284
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 8.056 46.758 8.256 ;
 END
 END vccd_1p0.gds284
 PIN vccd_1p0.gds285
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 8.0145 46.63 8.2145 ;
 END
 END vccd_1p0.gds285
 PIN vccd_1p0.gds286
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 10.244 50.33 10.444 ;
 END
 END vccd_1p0.gds286
 PIN vccd_1p0.gds287
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 8.984 50.33 9.184 ;
 END
 END vccd_1p0.gds287
 PIN vccd_1p0.gds288
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 7.724 50.33 7.924 ;
 END
 END vccd_1p0.gds288
 PIN vccd_1p0.gds289
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 6.464 50.33 6.664 ;
 END
 END vccd_1p0.gds289
 PIN vccd_1p0.gds290
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 8.0385 51.678 8.2385 ;
 END
 END vccd_1p0.gds290
 PIN vccd_1p0.gds291
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 8.0145 52.194 8.2145 ;
 END
 END vccd_1p0.gds291
 PIN vccd_1p0.gds292
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 8.056 52.066 8.256 ;
 END
 END vccd_1p0.gds292
 PIN vccd_1p0.gds293
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 7.9635 51.258 8.1635 ;
 END
 END vccd_1p0.gds293
 PIN vccd_1p0.gds294
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 8.06 51.838 8.26 ;
 END
 END vccd_1p0.gds294
 PIN vccd_1p0.gds295
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 8.0185 57.946 8.2185 ;
 END
 END vccd_1p0.gds295
 PIN vccd_1p0.gds296
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 6.4 65.134 6.6 ;
 END
 END vccd_1p0.gds296
 PIN vccd_1p0.gds297
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 10.18 65.134 10.38 ;
 END
 END vccd_1p0.gds297
 PIN vccd_1p0.gds298
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 8.92 65.134 9.12 ;
 END
 END vccd_1p0.gds298
 PIN vccd_1p0.gds299
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 7.66 65.134 7.86 ;
 END
 END vccd_1p0.gds299
 PIN vccd_1p0.gds300
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 7.86 64.894 8.06 ;
 END
 END vccd_1p0.gds300
 PIN vccd_1p0.gds301
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 7.9375 64.294 8.1375 ;
 END
 END vccd_1p0.gds301
 PIN vccd_1p0.gds302
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 8.06 64.054 8.26 ;
 END
 END vccd_1p0.gds302
 PIN vccd_1p0.gds303
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 8.056 63.81 8.256 ;
 END
 END vccd_1p0.gds303
 PIN vccd_1p0.gds304
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 8.0145 63.682 8.2145 ;
 END
 END vccd_1p0.gds304
 PIN vccd_1p0.gds305
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 10.244 67.382 10.444 ;
 END
 END vccd_1p0.gds305
 PIN vccd_1p0.gds306
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 10.18 65.554 10.38 ;
 END
 END vccd_1p0.gds306
 PIN vccd_1p0.gds307
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 10.3075 66.09 10.5075 ;
 END
 END vccd_1p0.gds307
 PIN vccd_1p0.gds308
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 8.984 67.382 9.184 ;
 END
 END vccd_1p0.gds308
 PIN vccd_1p0.gds309
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 8.92 65.554 9.12 ;
 END
 END vccd_1p0.gds309
 PIN vccd_1p0.gds310
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 9.0475 66.09 9.2475 ;
 END
 END vccd_1p0.gds310
 PIN vccd_1p0.gds311
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 7.724 67.382 7.924 ;
 END
 END vccd_1p0.gds311
 PIN vccd_1p0.gds312
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 7.66 65.554 7.86 ;
 END
 END vccd_1p0.gds312
 PIN vccd_1p0.gds313
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 7.7875 66.09 7.9875 ;
 END
 END vccd_1p0.gds313
 PIN vccd_1p0.gds314
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 6.464 67.382 6.664 ;
 END
 END vccd_1p0.gds314
 PIN vccd_1p0.gds315
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 6.4 65.554 6.6 ;
 END
 END vccd_1p0.gds315
 PIN vccd_1p0.gds316
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 6.5275 66.09 6.7275 ;
 END
 END vccd_1p0.gds316
 PIN vccd_1p0.gds317
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 8.112 66.446 8.312 ;
 END
 END vccd_1p0.gds317
 PIN vccd_1p0.gds318
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 8.112 65.898 8.312 ;
 END
 END vccd_1p0.gds318
 PIN vccd_1p0.gds319
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 8.0385 68.73 8.2385 ;
 END
 END vccd_1p0.gds319
 PIN vccd_1p0.gds320
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 8.0145 69.246 8.2145 ;
 END
 END vccd_1p0.gds320
 PIN vccd_1p0.gds321
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 8.056 69.118 8.256 ;
 END
 END vccd_1p0.gds321
 PIN vccd_1p0.gds322
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 7.9635 68.31 8.1635 ;
 END
 END vccd_1p0.gds322
 PIN vccd_1p0.gds323
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 8.094 66.898 8.294 ;
 END
 END vccd_1p0.gds323
 PIN vccd_1p0.gds324
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 8.094 66.654 8.294 ;
 END
 END vccd_1p0.gds324
 PIN vccd_1p0.gds325
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 8.06 68.89 8.26 ;
 END
 END vccd_1p0.gds325
 PIN vccd_1p0.gds326
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 13.058 0.43 13.258 ;
 END
 END vccd_1p0.gds326
 PIN vccd_1p0.gds327
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 14.873 1.542 15.073 ;
 END
 END vccd_1p0.gds327
 PIN vccd_1p0.gds328
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 14.7555 5.202 14.9555 ;
 END
 END vccd_1p0.gds328
 PIN vccd_1p0.gds329
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 13.613 1.542 13.813 ;
 END
 END vccd_1p0.gds329
 PIN vccd_1p0.gds330
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 13.4955 5.202 13.6955 ;
 END
 END vccd_1p0.gds330
 PIN vccd_1p0.gds331
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 12.353 1.542 12.553 ;
 END
 END vccd_1p0.gds331
 PIN vccd_1p0.gds332
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 12.2355 5.202 12.4355 ;
 END
 END vccd_1p0.gds332
 PIN vccd_1p0.gds333
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 11.093 1.542 11.293 ;
 END
 END vccd_1p0.gds333
 PIN vccd_1p0.gds334
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 10.9755 5.202 11.1755 ;
 END
 END vccd_1p0.gds334
 PIN vccd_1p0.gds335
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 13.169 0.548 13.369 ;
 END
 END vccd_1p0.gds335
 PIN vccd_1p0.gds336
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 13.1305 0.858 13.3305 ;
 END
 END vccd_1p0.gds336
 PIN vccd_1p0.gds337
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 12.968 1.362 13.168 ;
 END
 END vccd_1p0.gds337
 PIN vccd_1p0.gds338
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 13.186 1.782 13.386 ;
 END
 END vccd_1p0.gds338
 PIN vccd_1p0.gds339
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 13.067 1.218 13.267 ;
 END
 END vccd_1p0.gds339
 PIN vccd_1p0.gds340
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 13.141 1.962 13.341 ;
 END
 END vccd_1p0.gds340
 PIN vccd_1p0.gds341
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 13.0485 2.202 13.2485 ;
 END
 END vccd_1p0.gds341
 PIN vccd_1p0.gds342
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 13.1385 4.738 13.3385 ;
 END
 END vccd_1p0.gds342
 PIN vccd_1p0.gds343
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 13.0945 2.462 13.2945 ;
 END
 END vccd_1p0.gds343
 PIN vccd_1p0.gds344
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 13.087 2.622 13.287 ;
 END
 END vccd_1p0.gds344
 PIN vccd_1p0.gds345
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 13.087 1.09 13.287 ;
 END
 END vccd_1p0.gds345
 PIN vccd_1p0.gds346
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 12.9715 3.042 13.1715 ;
 END
 END vccd_1p0.gds346
 PIN vccd_1p0.gds347
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 13.1 2.882 13.3 ;
 END
 END vccd_1p0.gds347
 PIN vccd_1p0.gds348
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 13.06 3.39 13.26 ;
 END
 END vccd_1p0.gds348
 PIN vccd_1p0.gds349
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 13.096 3.262 13.296 ;
 END
 END vccd_1p0.gds349
 PIN vccd_1p0.gds350
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 13.139 3.666 13.339 ;
 END
 END vccd_1p0.gds350
 PIN vccd_1p0.gds351
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 13.1525 4.066 13.3525 ;
 END
 END vccd_1p0.gds351
 PIN vccd_1p0.gds352
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 13.1525 3.858 13.3525 ;
 END
 END vccd_1p0.gds352
 PIN vccd_1p0.gds353
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 13.1 4.258 13.3 ;
 END
 END vccd_1p0.gds353
 PIN vccd_1p0.gds354
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 13.138 4.546 13.338 ;
 END
 END vccd_1p0.gds354
 PIN vccd_1p0.gds355
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 13.162 5.01 13.362 ;
 END
 END vccd_1p0.gds355
 PIN vccd_1p0.gds356
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 4.34 11.308 4.396 11.508 ;
 RECT 4.76 11.284 4.816 11.484 ;
 RECT 5.096 11.308 5.152 11.508 ;
 RECT 4.34 12.568 4.396 12.768 ;
 RECT 4.76 12.544 4.816 12.744 ;
 RECT 5.096 12.568 5.152 12.768 ;
 RECT 4.34 13.828 4.396 14.028 ;
 RECT 4.76 13.804 4.816 14.004 ;
 RECT 5.096 13.828 5.152 14.028 ;
 RECT 4.34 15.088 4.396 15.288 ;
 RECT 4.76 15.064 4.816 15.264 ;
 RECT 5.096 15.088 5.152 15.288 ;
 RECT 3.584 14.8995 3.64 15.0995 ;
 RECT 4.172 14.9855 4.228 15.1855 ;
 RECT 4.928 14.942 4.984 15.142 ;
 RECT 3.584 13.6395 3.64 13.8395 ;
 RECT 4.172 13.7255 4.228 13.9255 ;
 RECT 4.928 13.682 4.984 13.882 ;
 RECT 3.584 12.3795 3.64 12.5795 ;
 RECT 4.172 12.4655 4.228 12.6655 ;
 RECT 4.928 12.422 4.984 12.622 ;
 RECT 3.584 11.1195 3.64 11.3195 ;
 RECT 4.172 11.2055 4.228 11.4055 ;
 RECT 4.928 11.162 4.984 11.362 ;
 END
 END vccd_1p0.gds356
 PIN vccd_1p0.gds357
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 13.1525 6.838 13.3525 ;
 END
 END vccd_1p0.gds357
 PIN vccd_1p0.gds358
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 13.162 6.05 13.362 ;
 END
 END vccd_1p0.gds358
 PIN vccd_1p0.gds359
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.754 13.1 5.794 13.3 ;
 END
 END vccd_1p0.gds359
 PIN vccd_1p0.gds360
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 13.189 6.306 13.389 ;
 END
 END vccd_1p0.gds360
 PIN vccd_1p0.gds361
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 13.1525 5.41 13.3525 ;
 END
 END vccd_1p0.gds361
 PIN vccd_1p0.gds362
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 13.1525 5.922 13.3525 ;
 END
 END vccd_1p0.gds362
 PIN vccd_1p0.gds363
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 13.042 5.602 13.242 ;
 END
 END vccd_1p0.gds363
 PIN vccd_1p0.gds364
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 13.079 6.582 13.279 ;
 END
 END vccd_1p0.gds364
 PIN vccd_1p0.gds365
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.6 14.9855 5.656 15.1855 ;
 RECT 5.264 14.9855 5.32 15.1855 ;
 RECT 5.432 14.8995 5.488 15.0995 ;
 RECT 5.936 14.8995 5.992 15.0995 ;
 RECT 5.768 14.8995 5.824 15.0995 ;
 RECT 6.44 14.914 6.496 15.114 ;
 RECT 6.272 14.8995 6.328 15.0995 ;
 RECT 6.104 15.088 6.16 15.288 ;
 RECT 5.6 13.7255 5.656 13.9255 ;
 RECT 5.264 13.7255 5.32 13.9255 ;
 RECT 5.432 13.6395 5.488 13.8395 ;
 RECT 5.936 13.6395 5.992 13.8395 ;
 RECT 5.768 13.6395 5.824 13.8395 ;
 RECT 6.44 13.654 6.496 13.854 ;
 RECT 6.272 13.6395 6.328 13.8395 ;
 RECT 6.104 13.828 6.16 14.028 ;
 RECT 5.6 12.4655 5.656 12.6655 ;
 RECT 5.264 12.4655 5.32 12.6655 ;
 RECT 5.432 12.3795 5.488 12.5795 ;
 RECT 5.936 12.3795 5.992 12.5795 ;
 RECT 5.768 12.3795 5.824 12.5795 ;
 RECT 6.44 12.394 6.496 12.594 ;
 RECT 6.272 12.3795 6.328 12.5795 ;
 RECT 6.104 12.568 6.16 12.768 ;
 RECT 5.6 11.2055 5.656 11.4055 ;
 RECT 5.264 11.2055 5.32 11.4055 ;
 RECT 5.432 11.1195 5.488 11.3195 ;
 RECT 5.936 11.1195 5.992 11.3195 ;
 RECT 5.768 11.1195 5.824 11.3195 ;
 RECT 6.44 11.134 6.496 11.334 ;
 RECT 6.272 11.1195 6.328 11.3195 ;
 RECT 6.104 11.308 6.16 11.508 ;
 END
 END vccd_1p0.gds365
 PIN vccd_1p0.gds366
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 11.44 13.978 11.64 ;
 END
 END vccd_1p0.gds366
 PIN vccd_1p0.gds367
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 12.7 13.978 12.9 ;
 END
 END vccd_1p0.gds367
 PIN vccd_1p0.gds368
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 13.96 13.978 14.16 ;
 END
 END vccd_1p0.gds368
 PIN vccd_1p0.gds369
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 15.22 13.978 15.42 ;
 END
 END vccd_1p0.gds369
 PIN vccd_1p0.gds370
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 15.22 14.398 15.42 ;
 END
 END vccd_1p0.gds370
 PIN vccd_1p0.gds371
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 15.3475 14.934 15.5475 ;
 END
 END vccd_1p0.gds371
 PIN vccd_1p0.gds372
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 13.96 14.398 14.16 ;
 END
 END vccd_1p0.gds372
 PIN vccd_1p0.gds373
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 14.0875 14.934 14.2875 ;
 END
 END vccd_1p0.gds373
 PIN vccd_1p0.gds374
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 12.7 14.398 12.9 ;
 END
 END vccd_1p0.gds374
 PIN vccd_1p0.gds375
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 12.8275 14.934 13.0275 ;
 END
 END vccd_1p0.gds375
 PIN vccd_1p0.gds376
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 11.44 14.398 11.64 ;
 END
 END vccd_1p0.gds376
 PIN vccd_1p0.gds377
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 11.5675 14.934 11.7675 ;
 END
 END vccd_1p0.gds377
 PIN vccd_1p0.gds378
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 13.152 14.742 13.352 ;
 END
 END vccd_1p0.gds378
 PIN vccd_1p0.gds379
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 12.9 13.738 13.1 ;
 END
 END vccd_1p0.gds379
 PIN vccd_1p0.gds380
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 13.1 12.898 13.3 ;
 END
 END vccd_1p0.gds380
 PIN vccd_1p0.gds381
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 12.9775 13.138 13.1775 ;
 END
 END vccd_1p0.gds381
 PIN vccd_1p0.gds382
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 13.096 12.654 13.296 ;
 END
 END vccd_1p0.gds382
 PIN vccd_1p0.gds383
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 13.0545 12.526 13.2545 ;
 END
 END vccd_1p0.gds383
 PIN vccd_1p0.gds384
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 15.284 16.226 15.484 ;
 END
 END vccd_1p0.gds384
 PIN vccd_1p0.gds385
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 14.024 16.226 14.224 ;
 END
 END vccd_1p0.gds385
 PIN vccd_1p0.gds386
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 12.764 16.226 12.964 ;
 END
 END vccd_1p0.gds386
 PIN vccd_1p0.gds387
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 11.504 16.226 11.704 ;
 END
 END vccd_1p0.gds387
 PIN vccd_1p0.gds388
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 13.134 15.742 13.334 ;
 END
 END vccd_1p0.gds388
 PIN vccd_1p0.gds389
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 13.152 15.29 13.352 ;
 END
 END vccd_1p0.gds389
 PIN vccd_1p0.gds390
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 13.0785 17.574 13.2785 ;
 END
 END vccd_1p0.gds390
 PIN vccd_1p0.gds391
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 13.0035 17.154 13.2035 ;
 END
 END vccd_1p0.gds391
 PIN vccd_1p0.gds392
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 13.1 17.734 13.3 ;
 END
 END vccd_1p0.gds392
 PIN vccd_1p0.gds393
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 13.134 15.498 13.334 ;
 END
 END vccd_1p0.gds393
 PIN vccd_1p0.gds394
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 13.096 17.962 13.296 ;
 END
 END vccd_1p0.gds394
 PIN vccd_1p0.gds395
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 13.0545 18.09 13.2545 ;
 END
 END vccd_1p0.gds395
 PIN vccd_1p0.gds396
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 13.0585 23.842 13.2585 ;
 END
 END vccd_1p0.gds396
 PIN vccd_1p0.gds397
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 13.1 29.95 13.3 ;
 END
 END vccd_1p0.gds397
 PIN vccd_1p0.gds398
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 13.096 29.706 13.296 ;
 END
 END vccd_1p0.gds398
 PIN vccd_1p0.gds399
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 13.0545 29.578 13.2545 ;
 END
 END vccd_1p0.gds399
 PIN vccd_1p0.gds400
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 15.22 31.03 15.42 ;
 END
 END vccd_1p0.gds400
 PIN vccd_1p0.gds401
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 13.96 31.03 14.16 ;
 END
 END vccd_1p0.gds401
 PIN vccd_1p0.gds402
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 12.7 31.03 12.9 ;
 END
 END vccd_1p0.gds402
 PIN vccd_1p0.gds403
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 11.44 31.03 11.64 ;
 END
 END vccd_1p0.gds403
 PIN vccd_1p0.gds404
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 11.504 33.278 11.704 ;
 END
 END vccd_1p0.gds404
 PIN vccd_1p0.gds405
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 11.44 31.45 11.64 ;
 END
 END vccd_1p0.gds405
 PIN vccd_1p0.gds406
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 11.5675 31.986 11.7675 ;
 END
 END vccd_1p0.gds406
 PIN vccd_1p0.gds407
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 12.764 33.278 12.964 ;
 END
 END vccd_1p0.gds407
 PIN vccd_1p0.gds408
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 12.7 31.45 12.9 ;
 END
 END vccd_1p0.gds408
 PIN vccd_1p0.gds409
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 12.8275 31.986 13.0275 ;
 END
 END vccd_1p0.gds409
 PIN vccd_1p0.gds410
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 14.024 33.278 14.224 ;
 END
 END vccd_1p0.gds410
 PIN vccd_1p0.gds411
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 13.96 31.45 14.16 ;
 END
 END vccd_1p0.gds411
 PIN vccd_1p0.gds412
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 14.0875 31.986 14.2875 ;
 END
 END vccd_1p0.gds412
 PIN vccd_1p0.gds413
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 15.284 33.278 15.484 ;
 END
 END vccd_1p0.gds413
 PIN vccd_1p0.gds414
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 15.22 31.45 15.42 ;
 END
 END vccd_1p0.gds414
 PIN vccd_1p0.gds415
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 15.3475 31.986 15.5475 ;
 END
 END vccd_1p0.gds415
 PIN vccd_1p0.gds416
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 12.9 30.79 13.1 ;
 END
 END vccd_1p0.gds416
 PIN vccd_1p0.gds417
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 12.9775 30.19 13.1775 ;
 END
 END vccd_1p0.gds417
 PIN vccd_1p0.gds418
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 13.152 32.342 13.352 ;
 END
 END vccd_1p0.gds418
 PIN vccd_1p0.gds419
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 13.152 31.794 13.352 ;
 END
 END vccd_1p0.gds419
 PIN vccd_1p0.gds420
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 13.0785 34.626 13.2785 ;
 END
 END vccd_1p0.gds420
 PIN vccd_1p0.gds421
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 13.0545 35.142 13.2545 ;
 END
 END vccd_1p0.gds421
 PIN vccd_1p0.gds422
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 13.096 35.014 13.296 ;
 END
 END vccd_1p0.gds422
 PIN vccd_1p0.gds423
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 13.0035 34.206 13.2035 ;
 END
 END vccd_1p0.gds423
 PIN vccd_1p0.gds424
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 13.134 32.794 13.334 ;
 END
 END vccd_1p0.gds424
 PIN vccd_1p0.gds425
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 13.134 32.55 13.334 ;
 END
 END vccd_1p0.gds425
 PIN vccd_1p0.gds426
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 13.1 34.786 13.3 ;
 END
 END vccd_1p0.gds426
 PIN vccd_1p0.gds427
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 13.0585 40.894 13.2585 ;
 END
 END vccd_1p0.gds427
 PIN vccd_1p0.gds428
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 11.44 48.082 11.64 ;
 END
 END vccd_1p0.gds428
 PIN vccd_1p0.gds429
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 12.7 48.082 12.9 ;
 END
 END vccd_1p0.gds429
 PIN vccd_1p0.gds430
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 13.96 48.082 14.16 ;
 END
 END vccd_1p0.gds430
 PIN vccd_1p0.gds431
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 15.22 48.502 15.42 ;
 END
 END vccd_1p0.gds431
 PIN vccd_1p0.gds432
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 15.3475 49.038 15.5475 ;
 END
 END vccd_1p0.gds432
 PIN vccd_1p0.gds433
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 13.96 48.502 14.16 ;
 END
 END vccd_1p0.gds433
 PIN vccd_1p0.gds434
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 14.0875 49.038 14.2875 ;
 END
 END vccd_1p0.gds434
 PIN vccd_1p0.gds435
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 12.7 48.502 12.9 ;
 END
 END vccd_1p0.gds435
 PIN vccd_1p0.gds436
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 12.8275 49.038 13.0275 ;
 END
 END vccd_1p0.gds436
 PIN vccd_1p0.gds437
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 11.44 48.502 11.64 ;
 END
 END vccd_1p0.gds437
 PIN vccd_1p0.gds438
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 11.5675 49.038 11.7675 ;
 END
 END vccd_1p0.gds438
 PIN vccd_1p0.gds439
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 15.22 48.082 15.42 ;
 END
 END vccd_1p0.gds439
 PIN vccd_1p0.gds440
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 12.9 47.842 13.1 ;
 END
 END vccd_1p0.gds440
 PIN vccd_1p0.gds441
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 12.9775 47.242 13.1775 ;
 END
 END vccd_1p0.gds441
 PIN vccd_1p0.gds442
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 13.152 49.394 13.352 ;
 END
 END vccd_1p0.gds442
 PIN vccd_1p0.gds443
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 13.152 48.846 13.352 ;
 END
 END vccd_1p0.gds443
 PIN vccd_1p0.gds444
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 13.134 49.846 13.334 ;
 END
 END vccd_1p0.gds444
 PIN vccd_1p0.gds445
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 13.134 49.602 13.334 ;
 END
 END vccd_1p0.gds445
 PIN vccd_1p0.gds446
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 13.1 47.002 13.3 ;
 END
 END vccd_1p0.gds446
 PIN vccd_1p0.gds447
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 13.096 46.758 13.296 ;
 END
 END vccd_1p0.gds447
 PIN vccd_1p0.gds448
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 13.0545 46.63 13.2545 ;
 END
 END vccd_1p0.gds448
 PIN vccd_1p0.gds449
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 15.284 50.33 15.484 ;
 END
 END vccd_1p0.gds449
 PIN vccd_1p0.gds450
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 14.024 50.33 14.224 ;
 END
 END vccd_1p0.gds450
 PIN vccd_1p0.gds451
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 12.764 50.33 12.964 ;
 END
 END vccd_1p0.gds451
 PIN vccd_1p0.gds452
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 11.504 50.33 11.704 ;
 END
 END vccd_1p0.gds452
 PIN vccd_1p0.gds453
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 13.0785 51.678 13.2785 ;
 END
 END vccd_1p0.gds453
 PIN vccd_1p0.gds454
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 13.0545 52.194 13.2545 ;
 END
 END vccd_1p0.gds454
 PIN vccd_1p0.gds455
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 13.096 52.066 13.296 ;
 END
 END vccd_1p0.gds455
 PIN vccd_1p0.gds456
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 13.0035 51.258 13.2035 ;
 END
 END vccd_1p0.gds456
 PIN vccd_1p0.gds457
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 13.1 51.838 13.3 ;
 END
 END vccd_1p0.gds457
 PIN vccd_1p0.gds458
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 13.0585 57.946 13.2585 ;
 END
 END vccd_1p0.gds458
 PIN vccd_1p0.gds459
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 15.22 65.134 15.42 ;
 END
 END vccd_1p0.gds459
 PIN vccd_1p0.gds460
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 13.96 65.134 14.16 ;
 END
 END vccd_1p0.gds460
 PIN vccd_1p0.gds461
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 12.7 65.134 12.9 ;
 END
 END vccd_1p0.gds461
 PIN vccd_1p0.gds462
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 11.44 65.134 11.64 ;
 END
 END vccd_1p0.gds462
 PIN vccd_1p0.gds463
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 12.9 64.894 13.1 ;
 END
 END vccd_1p0.gds463
 PIN vccd_1p0.gds464
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 12.9775 64.294 13.1775 ;
 END
 END vccd_1p0.gds464
 PIN vccd_1p0.gds465
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 13.1 64.054 13.3 ;
 END
 END vccd_1p0.gds465
 PIN vccd_1p0.gds466
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 13.096 63.81 13.296 ;
 END
 END vccd_1p0.gds466
 PIN vccd_1p0.gds467
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 13.0545 63.682 13.2545 ;
 END
 END vccd_1p0.gds467
 PIN vccd_1p0.gds468
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 15.284 67.382 15.484 ;
 END
 END vccd_1p0.gds468
 PIN vccd_1p0.gds469
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 15.22 65.554 15.42 ;
 END
 END vccd_1p0.gds469
 PIN vccd_1p0.gds470
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 15.3475 66.09 15.5475 ;
 END
 END vccd_1p0.gds470
 PIN vccd_1p0.gds471
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 14.024 67.382 14.224 ;
 END
 END vccd_1p0.gds471
 PIN vccd_1p0.gds472
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 13.96 65.554 14.16 ;
 END
 END vccd_1p0.gds472
 PIN vccd_1p0.gds473
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 14.0875 66.09 14.2875 ;
 END
 END vccd_1p0.gds473
 PIN vccd_1p0.gds474
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 12.764 67.382 12.964 ;
 END
 END vccd_1p0.gds474
 PIN vccd_1p0.gds475
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 12.7 65.554 12.9 ;
 END
 END vccd_1p0.gds475
 PIN vccd_1p0.gds476
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 12.8275 66.09 13.0275 ;
 END
 END vccd_1p0.gds476
 PIN vccd_1p0.gds477
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 11.504 67.382 11.704 ;
 END
 END vccd_1p0.gds477
 PIN vccd_1p0.gds478
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 11.44 65.554 11.64 ;
 END
 END vccd_1p0.gds478
 PIN vccd_1p0.gds479
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 11.5675 66.09 11.7675 ;
 END
 END vccd_1p0.gds479
 PIN vccd_1p0.gds480
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 13.152 66.446 13.352 ;
 END
 END vccd_1p0.gds480
 PIN vccd_1p0.gds481
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 13.152 65.898 13.352 ;
 END
 END vccd_1p0.gds481
 PIN vccd_1p0.gds482
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 13.0785 68.73 13.2785 ;
 END
 END vccd_1p0.gds482
 PIN vccd_1p0.gds483
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 13.0545 69.246 13.2545 ;
 END
 END vccd_1p0.gds483
 PIN vccd_1p0.gds484
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 13.096 69.118 13.296 ;
 END
 END vccd_1p0.gds484
 PIN vccd_1p0.gds485
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 13.0035 68.31 13.2035 ;
 END
 END vccd_1p0.gds485
 PIN vccd_1p0.gds486
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 13.134 66.898 13.334 ;
 END
 END vccd_1p0.gds486
 PIN vccd_1p0.gds487
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 13.134 66.654 13.334 ;
 END
 END vccd_1p0.gds487
 PIN vccd_1p0.gds488
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 13.1 68.89 13.3 ;
 END
 END vccd_1p0.gds488
 PIN vccd_1p0.gds489
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 18.098 0.43 18.298 ;
 END
 END vccd_1p0.gds489
 PIN vccd_1p0.gds490
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 19.913 1.542 20.113 ;
 END
 END vccd_1p0.gds490
 PIN vccd_1p0.gds491
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 16.133 1.542 16.333 ;
 END
 END vccd_1p0.gds491
 PIN vccd_1p0.gds492
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 16.0155 5.202 16.2155 ;
 END
 END vccd_1p0.gds492
 PIN vccd_1p0.gds493
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 17.393 1.542 17.593 ;
 END
 END vccd_1p0.gds493
 PIN vccd_1p0.gds494
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 17.2755 5.202 17.4755 ;
 END
 END vccd_1p0.gds494
 PIN vccd_1p0.gds495
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 18.653 1.542 18.853 ;
 END
 END vccd_1p0.gds495
 PIN vccd_1p0.gds496
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 18.5355 5.202 18.7355 ;
 END
 END vccd_1p0.gds496
 PIN vccd_1p0.gds497
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 18.3535 0.548 18.5535 ;
 END
 END vccd_1p0.gds497
 PIN vccd_1p0.gds498
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 18.1705 0.858 18.3705 ;
 END
 END vccd_1p0.gds498
 PIN vccd_1p0.gds499
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 18.008 1.362 18.208 ;
 END
 END vccd_1p0.gds499
 PIN vccd_1p0.gds500
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 18.342 1.782 18.542 ;
 END
 END vccd_1p0.gds500
 PIN vccd_1p0.gds501
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 18.107 1.218 18.307 ;
 END
 END vccd_1p0.gds501
 PIN vccd_1p0.gds502
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 18.181 1.962 18.381 ;
 END
 END vccd_1p0.gds502
 PIN vccd_1p0.gds503
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 18.0885 2.202 18.2885 ;
 END
 END vccd_1p0.gds503
 PIN vccd_1p0.gds504
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 19.885 5.202 20.085 ;
 END
 END vccd_1p0.gds504
 PIN vccd_1p0.gds505
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 18.1785 4.738 18.3785 ;
 END
 END vccd_1p0.gds505
 PIN vccd_1p0.gds506
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 18.1345 2.462 18.3345 ;
 END
 END vccd_1p0.gds506
 PIN vccd_1p0.gds507
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 18.127 2.622 18.327 ;
 END
 END vccd_1p0.gds507
 PIN vccd_1p0.gds508
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 18.127 1.09 18.327 ;
 END
 END vccd_1p0.gds508
 PIN vccd_1p0.gds509
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 18.0115 3.042 18.2115 ;
 END
 END vccd_1p0.gds509
 PIN vccd_1p0.gds510
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 18.14 2.882 18.34 ;
 END
 END vccd_1p0.gds510
 PIN vccd_1p0.gds511
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 18.1 3.39 18.3 ;
 END
 END vccd_1p0.gds511
 PIN vccd_1p0.gds512
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 18.136 3.262 18.336 ;
 END
 END vccd_1p0.gds512
 PIN vccd_1p0.gds513
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 18.179 3.666 18.379 ;
 END
 END vccd_1p0.gds513
 PIN vccd_1p0.gds514
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 18.1925 4.066 18.3925 ;
 END
 END vccd_1p0.gds514
 PIN vccd_1p0.gds515
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 18.1925 3.858 18.3925 ;
 END
 END vccd_1p0.gds515
 PIN vccd_1p0.gds516
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 18.14 4.258 18.34 ;
 END
 END vccd_1p0.gds516
 PIN vccd_1p0.gds517
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 18.178 4.546 18.378 ;
 END
 END vccd_1p0.gds517
 PIN vccd_1p0.gds518
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 18.202 5.01 18.402 ;
 END
 END vccd_1p0.gds518
 PIN vccd_1p0.gds519
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 4.34 16.348 4.396 16.548 ;
 RECT 4.76 16.324 4.816 16.524 ;
 RECT 5.096 16.348 5.152 16.548 ;
 RECT 4.34 17.608 4.396 17.808 ;
 RECT 4.76 17.584 4.816 17.784 ;
 RECT 5.096 17.608 5.152 17.808 ;
 RECT 4.34 18.868 4.396 19.068 ;
 RECT 4.76 18.844 4.816 19.044 ;
 RECT 5.096 18.868 5.152 19.068 ;
 RECT 4.34 20.128 4.396 20.328 ;
 RECT 4.76 20.104 4.816 20.304 ;
 RECT 5.096 20.128 5.152 20.328 ;
 RECT 3.584 19.9395 3.64 20.1395 ;
 RECT 4.172 20.0255 4.228 20.2255 ;
 RECT 4.928 19.982 4.984 20.182 ;
 RECT 3.584 18.6795 3.64 18.8795 ;
 RECT 4.172 18.7655 4.228 18.9655 ;
 RECT 4.928 18.722 4.984 18.922 ;
 RECT 3.584 17.4195 3.64 17.6195 ;
 RECT 4.172 17.5055 4.228 17.7055 ;
 RECT 4.928 17.462 4.984 17.662 ;
 RECT 3.584 16.1595 3.64 16.3595 ;
 RECT 4.172 16.2455 4.228 16.4455 ;
 RECT 4.928 16.202 4.984 16.402 ;
 END
 END vccd_1p0.gds519
 PIN vccd_1p0.gds520
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 18.1925 6.838 18.3925 ;
 END
 END vccd_1p0.gds520
 PIN vccd_1p0.gds521
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 18.202 6.05 18.402 ;
 END
 END vccd_1p0.gds521
 PIN vccd_1p0.gds522
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.754 18.14 5.794 18.34 ;
 END
 END vccd_1p0.gds522
 PIN vccd_1p0.gds523
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 18.229 6.306 18.429 ;
 END
 END vccd_1p0.gds523
 PIN vccd_1p0.gds524
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 18.1925 5.41 18.3925 ;
 END
 END vccd_1p0.gds524
 PIN vccd_1p0.gds525
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 18.1925 5.922 18.3925 ;
 END
 END vccd_1p0.gds525
 PIN vccd_1p0.gds526
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 18.082 5.602 18.282 ;
 END
 END vccd_1p0.gds526
 PIN vccd_1p0.gds527
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 18.119 6.582 18.319 ;
 END
 END vccd_1p0.gds527
 PIN vccd_1p0.gds528
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.6 20.0255 5.656 20.2255 ;
 RECT 5.264 20.0255 5.32 20.2255 ;
 RECT 5.432 19.9395 5.488 20.1395 ;
 RECT 5.936 19.9395 5.992 20.1395 ;
 RECT 5.768 19.9395 5.824 20.1395 ;
 RECT 6.44 19.954 6.496 20.154 ;
 RECT 6.272 19.9395 6.328 20.1395 ;
 RECT 6.104 20.128 6.16 20.328 ;
 RECT 5.6 18.7655 5.656 18.9655 ;
 RECT 5.264 18.7655 5.32 18.9655 ;
 RECT 5.432 18.6795 5.488 18.8795 ;
 RECT 5.936 18.6795 5.992 18.8795 ;
 RECT 5.768 18.6795 5.824 18.8795 ;
 RECT 6.44 18.694 6.496 18.894 ;
 RECT 6.272 18.6795 6.328 18.8795 ;
 RECT 6.104 18.868 6.16 19.068 ;
 RECT 5.6 17.5055 5.656 17.7055 ;
 RECT 5.264 17.5055 5.32 17.7055 ;
 RECT 5.432 17.4195 5.488 17.6195 ;
 RECT 5.936 17.4195 5.992 17.6195 ;
 RECT 5.768 17.4195 5.824 17.6195 ;
 RECT 6.44 17.434 6.496 17.634 ;
 RECT 6.272 17.4195 6.328 17.6195 ;
 RECT 6.104 17.608 6.16 17.808 ;
 RECT 5.6 16.2455 5.656 16.4455 ;
 RECT 5.264 16.2455 5.32 16.4455 ;
 RECT 5.432 16.1595 5.488 16.3595 ;
 RECT 5.936 16.1595 5.992 16.3595 ;
 RECT 5.768 16.1595 5.824 16.3595 ;
 RECT 6.44 16.174 6.496 16.374 ;
 RECT 6.272 16.1595 6.328 16.3595 ;
 RECT 6.104 16.348 6.16 16.548 ;
 END
 END vccd_1p0.gds528
 PIN vccd_1p0.gds529
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 19 13.978 19.2 ;
 END
 END vccd_1p0.gds529
 PIN vccd_1p0.gds530
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 20.26 13.978 20.46 ;
 END
 END vccd_1p0.gds530
 PIN vccd_1p0.gds531
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 19 14.398 19.2 ;
 END
 END vccd_1p0.gds531
 PIN vccd_1p0.gds532
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 20.3805 14.398 20.5805 ;
 END
 END vccd_1p0.gds532
 PIN vccd_1p0.gds533
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 17.74 13.978 17.94 ;
 END
 END vccd_1p0.gds533
 PIN vccd_1p0.gds534
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 16.48 14.398 16.68 ;
 END
 END vccd_1p0.gds534
 PIN vccd_1p0.gds535
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 16.6075 14.934 16.8075 ;
 END
 END vccd_1p0.gds535
 PIN vccd_1p0.gds536
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 17.74 14.398 17.94 ;
 END
 END vccd_1p0.gds536
 PIN vccd_1p0.gds537
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 17.8675 14.934 18.0675 ;
 END
 END vccd_1p0.gds537
 PIN vccd_1p0.gds538
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 18.192 14.742 18.392 ;
 END
 END vccd_1p0.gds538
 PIN vccd_1p0.gds539
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 16.48 13.978 16.68 ;
 END
 END vccd_1p0.gds539
 PIN vccd_1p0.gds540
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 17.94 13.738 18.14 ;
 END
 END vccd_1p0.gds540
 PIN vccd_1p0.gds541
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 18.14 12.898 18.34 ;
 END
 END vccd_1p0.gds541
 PIN vccd_1p0.gds542
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 18.0175 13.138 18.2175 ;
 END
 END vccd_1p0.gds542
 PIN vccd_1p0.gds543
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 18.136 12.654 18.336 ;
 END
 END vccd_1p0.gds543
 PIN vccd_1p0.gds544
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 18.0945 12.526 18.2945 ;
 END
 END vccd_1p0.gds544
 PIN vccd_1p0.gds545
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 19.1275 14.934 19.3275 ;
 END
 END vccd_1p0.gds545
 PIN vccd_1p0.gds546
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 19.064 16.226 19.264 ;
 END
 END vccd_1p0.gds546
 PIN vccd_1p0.gds547
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 17.804 16.226 18.004 ;
 END
 END vccd_1p0.gds547
 PIN vccd_1p0.gds548
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 16.544 16.226 16.744 ;
 END
 END vccd_1p0.gds548
 PIN vccd_1p0.gds549
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 18.174 15.742 18.374 ;
 END
 END vccd_1p0.gds549
 PIN vccd_1p0.gds550
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 18.192 15.29 18.392 ;
 END
 END vccd_1p0.gds550
 PIN vccd_1p0.gds551
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 18.1185 17.574 18.3185 ;
 END
 END vccd_1p0.gds551
 PIN vccd_1p0.gds552
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 18.0435 17.154 18.2435 ;
 END
 END vccd_1p0.gds552
 PIN vccd_1p0.gds553
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 18.14 17.734 18.34 ;
 END
 END vccd_1p0.gds553
 PIN vccd_1p0.gds554
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 18.174 15.498 18.374 ;
 END
 END vccd_1p0.gds554
 PIN vccd_1p0.gds555
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 18.136 17.962 18.336 ;
 END
 END vccd_1p0.gds555
 PIN vccd_1p0.gds556
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 18.0945 18.09 18.2945 ;
 END
 END vccd_1p0.gds556
 PIN vccd_1p0.gds557
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 18.0985 23.842 18.2985 ;
 END
 END vccd_1p0.gds557
 PIN vccd_1p0.gds558
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 18.14 29.95 18.34 ;
 END
 END vccd_1p0.gds558
 PIN vccd_1p0.gds559
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 18.136 29.706 18.336 ;
 END
 END vccd_1p0.gds559
 PIN vccd_1p0.gds560
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 18.0945 29.578 18.2945 ;
 END
 END vccd_1p0.gds560
 PIN vccd_1p0.gds561
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 19 31.03 19.2 ;
 END
 END vccd_1p0.gds561
 PIN vccd_1p0.gds562
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 20.26 31.03 20.46 ;
 END
 END vccd_1p0.gds562
 PIN vccd_1p0.gds563
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 19.064 33.278 19.264 ;
 END
 END vccd_1p0.gds563
 PIN vccd_1p0.gds564
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 19 31.45 19.2 ;
 END
 END vccd_1p0.gds564
 PIN vccd_1p0.gds565
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 17.74 31.03 17.94 ;
 END
 END vccd_1p0.gds565
 PIN vccd_1p0.gds566
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 16.48 31.03 16.68 ;
 END
 END vccd_1p0.gds566
 PIN vccd_1p0.gds567
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 16.544 33.278 16.744 ;
 END
 END vccd_1p0.gds567
 PIN vccd_1p0.gds568
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 16.48 31.45 16.68 ;
 END
 END vccd_1p0.gds568
 PIN vccd_1p0.gds569
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 16.6075 31.986 16.8075 ;
 END
 END vccd_1p0.gds569
 PIN vccd_1p0.gds570
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 17.804 33.278 18.004 ;
 END
 END vccd_1p0.gds570
 PIN vccd_1p0.gds571
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 17.74 31.45 17.94 ;
 END
 END vccd_1p0.gds571
 PIN vccd_1p0.gds572
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 17.8675 31.986 18.0675 ;
 END
 END vccd_1p0.gds572
 PIN vccd_1p0.gds573
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 17.94 30.79 18.14 ;
 END
 END vccd_1p0.gds573
 PIN vccd_1p0.gds574
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 18.0175 30.19 18.2175 ;
 END
 END vccd_1p0.gds574
 PIN vccd_1p0.gds575
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 18.192 32.342 18.392 ;
 END
 END vccd_1p0.gds575
 PIN vccd_1p0.gds576
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 20.3805 31.45 20.5805 ;
 END
 END vccd_1p0.gds576
 PIN vccd_1p0.gds577
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 18.192 31.794 18.392 ;
 END
 END vccd_1p0.gds577
 PIN vccd_1p0.gds578
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 18.1185 34.626 18.3185 ;
 END
 END vccd_1p0.gds578
 PIN vccd_1p0.gds579
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 18.0945 35.142 18.2945 ;
 END
 END vccd_1p0.gds579
 PIN vccd_1p0.gds580
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 19.1275 31.986 19.3275 ;
 END
 END vccd_1p0.gds580
 PIN vccd_1p0.gds581
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 18.136 35.014 18.336 ;
 END
 END vccd_1p0.gds581
 PIN vccd_1p0.gds582
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 18.0435 34.206 18.2435 ;
 END
 END vccd_1p0.gds582
 PIN vccd_1p0.gds583
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 18.174 32.794 18.374 ;
 END
 END vccd_1p0.gds583
 PIN vccd_1p0.gds584
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 18.174 32.55 18.374 ;
 END
 END vccd_1p0.gds584
 PIN vccd_1p0.gds585
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 18.14 34.786 18.34 ;
 END
 END vccd_1p0.gds585
 PIN vccd_1p0.gds586
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 18.0985 40.894 18.2985 ;
 END
 END vccd_1p0.gds586
 PIN vccd_1p0.gds587
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 19 48.082 19.2 ;
 END
 END vccd_1p0.gds587
 PIN vccd_1p0.gds588
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 20.26 48.082 20.46 ;
 END
 END vccd_1p0.gds588
 PIN vccd_1p0.gds589
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 19 48.502 19.2 ;
 END
 END vccd_1p0.gds589
 PIN vccd_1p0.gds590
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 17.74 48.082 17.94 ;
 END
 END vccd_1p0.gds590
 PIN vccd_1p0.gds591
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 16.48 48.502 16.68 ;
 END
 END vccd_1p0.gds591
 PIN vccd_1p0.gds592
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 16.6075 49.038 16.8075 ;
 END
 END vccd_1p0.gds592
 PIN vccd_1p0.gds593
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 17.74 48.502 17.94 ;
 END
 END vccd_1p0.gds593
 PIN vccd_1p0.gds594
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 17.8675 49.038 18.0675 ;
 END
 END vccd_1p0.gds594
 PIN vccd_1p0.gds595
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 16.48 48.082 16.68 ;
 END
 END vccd_1p0.gds595
 PIN vccd_1p0.gds596
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 17.94 47.842 18.14 ;
 END
 END vccd_1p0.gds596
 PIN vccd_1p0.gds597
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 18.0175 47.242 18.2175 ;
 END
 END vccd_1p0.gds597
 PIN vccd_1p0.gds598
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 18.192 49.394 18.392 ;
 END
 END vccd_1p0.gds598
 PIN vccd_1p0.gds599
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 20.3805 48.502 20.5805 ;
 END
 END vccd_1p0.gds599
 PIN vccd_1p0.gds600
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 18.192 48.846 18.392 ;
 END
 END vccd_1p0.gds600
 PIN vccd_1p0.gds601
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 19.1275 49.038 19.3275 ;
 END
 END vccd_1p0.gds601
 PIN vccd_1p0.gds602
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 18.174 49.846 18.374 ;
 END
 END vccd_1p0.gds602
 PIN vccd_1p0.gds603
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 18.174 49.602 18.374 ;
 END
 END vccd_1p0.gds603
 PIN vccd_1p0.gds604
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 18.14 47.002 18.34 ;
 END
 END vccd_1p0.gds604
 PIN vccd_1p0.gds605
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 18.136 46.758 18.336 ;
 END
 END vccd_1p0.gds605
 PIN vccd_1p0.gds606
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 18.0945 46.63 18.2945 ;
 END
 END vccd_1p0.gds606
 PIN vccd_1p0.gds607
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 19.064 50.33 19.264 ;
 END
 END vccd_1p0.gds607
 PIN vccd_1p0.gds608
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 16.544 50.33 16.744 ;
 END
 END vccd_1p0.gds608
 PIN vccd_1p0.gds609
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 17.804 50.33 18.004 ;
 END
 END vccd_1p0.gds609
 PIN vccd_1p0.gds610
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 18.1185 51.678 18.3185 ;
 END
 END vccd_1p0.gds610
 PIN vccd_1p0.gds611
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 18.0945 52.194 18.2945 ;
 END
 END vccd_1p0.gds611
 PIN vccd_1p0.gds612
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 18.136 52.066 18.336 ;
 END
 END vccd_1p0.gds612
 PIN vccd_1p0.gds613
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 18.0435 51.258 18.2435 ;
 END
 END vccd_1p0.gds613
 PIN vccd_1p0.gds614
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 18.14 51.838 18.34 ;
 END
 END vccd_1p0.gds614
 PIN vccd_1p0.gds615
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 18.0985 57.946 18.2985 ;
 END
 END vccd_1p0.gds615
 PIN vccd_1p0.gds616
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 19 65.134 19.2 ;
 END
 END vccd_1p0.gds616
 PIN vccd_1p0.gds617
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 20.26 65.134 20.46 ;
 END
 END vccd_1p0.gds617
 PIN vccd_1p0.gds618
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 17.74 65.134 17.94 ;
 END
 END vccd_1p0.gds618
 PIN vccd_1p0.gds619
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 16.48 65.134 16.68 ;
 END
 END vccd_1p0.gds619
 PIN vccd_1p0.gds620
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 17.94 64.894 18.14 ;
 END
 END vccd_1p0.gds620
 PIN vccd_1p0.gds621
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 18.0175 64.294 18.2175 ;
 END
 END vccd_1p0.gds621
 PIN vccd_1p0.gds622
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 18.14 64.054 18.34 ;
 END
 END vccd_1p0.gds622
 PIN vccd_1p0.gds623
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 18.136 63.81 18.336 ;
 END
 END vccd_1p0.gds623
 PIN vccd_1p0.gds624
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 18.0945 63.682 18.2945 ;
 END
 END vccd_1p0.gds624
 PIN vccd_1p0.gds625
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 19.064 67.382 19.264 ;
 END
 END vccd_1p0.gds625
 PIN vccd_1p0.gds626
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 19 65.554 19.2 ;
 END
 END vccd_1p0.gds626
 PIN vccd_1p0.gds627
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 17.804 67.382 18.004 ;
 END
 END vccd_1p0.gds627
 PIN vccd_1p0.gds628
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 17.74 65.554 17.94 ;
 END
 END vccd_1p0.gds628
 PIN vccd_1p0.gds629
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 17.8675 66.09 18.0675 ;
 END
 END vccd_1p0.gds629
 PIN vccd_1p0.gds630
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 16.544 67.382 16.744 ;
 END
 END vccd_1p0.gds630
 PIN vccd_1p0.gds631
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 16.48 65.554 16.68 ;
 END
 END vccd_1p0.gds631
 PIN vccd_1p0.gds632
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 16.6075 66.09 16.8075 ;
 END
 END vccd_1p0.gds632
 PIN vccd_1p0.gds633
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 18.192 66.446 18.392 ;
 END
 END vccd_1p0.gds633
 PIN vccd_1p0.gds634
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 20.3805 65.554 20.5805 ;
 END
 END vccd_1p0.gds634
 PIN vccd_1p0.gds635
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 18.192 65.898 18.392 ;
 END
 END vccd_1p0.gds635
 PIN vccd_1p0.gds636
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 18.1185 68.73 18.3185 ;
 END
 END vccd_1p0.gds636
 PIN vccd_1p0.gds637
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 18.0945 69.246 18.2945 ;
 END
 END vccd_1p0.gds637
 PIN vccd_1p0.gds638
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 19.1275 66.09 19.3275 ;
 END
 END vccd_1p0.gds638
 PIN vccd_1p0.gds639
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 18.136 69.118 18.336 ;
 END
 END vccd_1p0.gds639
 PIN vccd_1p0.gds640
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 18.0435 68.31 18.2435 ;
 END
 END vccd_1p0.gds640
 PIN vccd_1p0.gds641
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 18.174 66.898 18.374 ;
 END
 END vccd_1p0.gds641
 PIN vccd_1p0.gds642
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 18.174 66.654 18.374 ;
 END
 END vccd_1p0.gds642
 PIN vccd_1p0.gds643
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 18.14 68.89 18.34 ;
 END
 END vccd_1p0.gds643
 PIN vccd_1p0.gds644
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 23.749 0.43 23.949 ;
 END
 END vccd_1p0.gds644
 PIN vccd_1p0.gds645
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 23.444 0.548 23.644 ;
 END
 END vccd_1p0.gds645
 PIN vccd_1p0.gds646
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 23.18 1.542 23.38 ;
 END
 END vccd_1p0.gds646
 PIN vccd_1p0.gds647
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 23.112 0.858 23.312 ;
 END
 END vccd_1p0.gds647
 PIN vccd_1p0.gds648
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 23.177 1.362 23.377 ;
 END
 END vccd_1p0.gds648
 PIN vccd_1p0.gds649
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 21.09 1.782 21.29 ;
 END
 END vccd_1p0.gds649
 PIN vccd_1p0.gds650
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 23.2035 1.218 23.4035 ;
 END
 END vccd_1p0.gds650
 PIN vccd_1p0.gds651
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 22.904 1.962 23.104 ;
 END
 END vccd_1p0.gds651
 PIN vccd_1p0.gds652
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 21.1605 4.738 21.3605 ;
 END
 END vccd_1p0.gds652
 PIN vccd_1p0.gds653
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 22.829 2.462 23.029 ;
 END
 END vccd_1p0.gds653
 PIN vccd_1p0.gds654
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 21.117 2.622 21.317 ;
 END
 END vccd_1p0.gds654
 PIN vccd_1p0.gds655
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 23.184 1.09 23.384 ;
 END
 END vccd_1p0.gds655
 PIN vccd_1p0.gds656
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 23.197 3.042 23.397 ;
 END
 END vccd_1p0.gds656
 PIN vccd_1p0.gds657
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 23.58 2.882 23.78 ;
 END
 END vccd_1p0.gds657
 PIN vccd_1p0.gds658
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 23.144 3.39 23.344 ;
 END
 END vccd_1p0.gds658
 PIN vccd_1p0.gds659
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 22.85 2.622 23.05 ;
 END
 END vccd_1p0.gds659
 PIN vccd_1p0.gds660
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 23.2815 3.262 23.4815 ;
 END
 END vccd_1p0.gds660
 PIN vccd_1p0.gds661
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 21.3375 3.666 21.5375 ;
 END
 END vccd_1p0.gds661
 PIN vccd_1p0.gds662
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 21.299 4.066 21.499 ;
 END
 END vccd_1p0.gds662
 PIN vccd_1p0.gds663
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 23.4305 3.858 23.6305 ;
 END
 END vccd_1p0.gds663
 PIN vccd_1p0.gds664
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 20.879 4.258 21.079 ;
 END
 END vccd_1p0.gds664
 PIN vccd_1p0.gds665
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 23.2685 4.546 23.4685 ;
 END
 END vccd_1p0.gds665
 PIN vccd_1p0.gds666
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 23.4755 5.01 23.6755 ;
 END
 END vccd_1p0.gds666
 PIN vccd_1p0.gds667
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.982 25.238 10.022 25.438 ;
 END
 END vccd_1p0.gds667
 PIN vccd_1p0.gds668
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.31 25.238 9.35 25.438 ;
 END
 END vccd_1p0.gds668
 PIN vccd_1p0.gds669
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.638 25.238 8.678 25.438 ;
 END
 END vccd_1p0.gds669
 PIN vccd_1p0.gds670
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.966 25.238 8.006 25.438 ;
 END
 END vccd_1p0.gds670
 PIN vccd_1p0.gds671
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.294 25.238 7.334 25.438 ;
 END
 END vccd_1p0.gds671
 PIN vccd_1p0.gds672
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.046 21.826 10.086 22.026 ;
 END
 END vccd_1p0.gds672
 PIN vccd_1p0.gds673
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.374 21.826 9.414 22.026 ;
 END
 END vccd_1p0.gds673
 PIN vccd_1p0.gds674
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.702 21.826 8.742 22.026 ;
 END
 END vccd_1p0.gds674
 PIN vccd_1p0.gds675
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.03 21.826 8.07 22.026 ;
 END
 END vccd_1p0.gds675
 PIN vccd_1p0.gds676
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.848 22.8795 9.894 23.0795 ;
 END
 END vccd_1p0.gds676
 PIN vccd_1p0.gds677
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.176 22.8795 9.222 23.0795 ;
 END
 END vccd_1p0.gds677
 PIN vccd_1p0.gds678
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.504 22.8795 8.55 23.0795 ;
 END
 END vccd_1p0.gds678
 PIN vccd_1p0.gds679
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.832 22.8795 7.878 23.0795 ;
 END
 END vccd_1p0.gds679
 PIN vccd_1p0.gds680
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.16 22.901 7.206 23.101 ;
 END
 END vccd_1p0.gds680
 PIN vccd_1p0.gds681
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 22.6595 6.838 22.8595 ;
 END
 END vccd_1p0.gds681
 PIN vccd_1p0.gds682
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 21.1485 6.05 21.3485 ;
 END
 END vccd_1p0.gds682
 PIN vccd_1p0.gds683
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 20.666 6.306 20.866 ;
 END
 END vccd_1p0.gds683
 PIN vccd_1p0.gds684
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 21.565 5.41 21.765 ;
 END
 END vccd_1p0.gds684
 PIN vccd_1p0.gds685
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 21.247 5.922 21.447 ;
 END
 END vccd_1p0.gds685
 PIN vccd_1p0.gds686
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 23.4065 5.602 23.6065 ;
 END
 END vccd_1p0.gds686
 PIN vccd_1p0.gds687
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 24.1075 6.306 24.3075 ;
 END
 END vccd_1p0.gds687
 PIN vccd_1p0.gds688
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.358 22.112 7.398 22.312 ;
 END
 END vccd_1p0.gds688
 PIN vccd_1p0.gds689
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 23.291 6.582 23.491 ;
 END
 END vccd_1p0.gds689
 PIN vccd_1p0.gds690
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.998 25.238 12.038 25.438 ;
 END
 END vccd_1p0.gds690
 PIN vccd_1p0.gds691
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.326 25.238 11.366 25.438 ;
 END
 END vccd_1p0.gds691
 PIN vccd_1p0.gds692
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.654 25.238 10.694 25.438 ;
 END
 END vccd_1p0.gds692
 PIN vccd_1p0.gds693
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.062 21.8735 12.102 22.0735 ;
 END
 END vccd_1p0.gds693
 PIN vccd_1p0.gds694
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.39 21.826 11.43 22.026 ;
 END
 END vccd_1p0.gds694
 PIN vccd_1p0.gds695
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.718 21.826 10.758 22.026 ;
 END
 END vccd_1p0.gds695
 PIN vccd_1p0.gds696
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 24.432 13.138 24.632 ;
 END
 END vccd_1p0.gds696
 PIN vccd_1p0.gds697
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 24.056 12.654 24.256 ;
 END
 END vccd_1p0.gds697
 PIN vccd_1p0.gds698
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 23.3505 15.29 23.5505 ;
 END
 END vccd_1p0.gds698
 PIN vccd_1p0.gds699
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 22.7035 14.934 22.9035 ;
 END
 END vccd_1p0.gds699
 PIN vccd_1p0.gds700
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.678 22.434 12.718 22.634 ;
 END
 END vccd_1p0.gds700
 PIN vccd_1p0.gds701
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.262 21.013 13.318 21.213 ;
 END
 END vccd_1p0.gds701
 PIN vccd_1p0.gds702
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 21.573 13.978 21.773 ;
 END
 END vccd_1p0.gds702
 PIN vccd_1p0.gds703
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 20.9785 14.742 21.1785 ;
 END
 END vccd_1p0.gds703
 PIN vccd_1p0.gds704
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 20.738 13.738 20.938 ;
 END
 END vccd_1p0.gds704
 PIN vccd_1p0.gds705
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 20.984 12.898 21.184 ;
 END
 END vccd_1p0.gds705
 PIN vccd_1p0.gds706
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 20.737 12.526 20.937 ;
 END
 END vccd_1p0.gds706
 PIN vccd_1p0.gds707
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 20.5055 14.934 20.7055 ;
 END
 END vccd_1p0.gds707
 PIN vccd_1p0.gds708
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.864 22.8795 11.91 23.0795 ;
 END
 END vccd_1p0.gds708
 PIN vccd_1p0.gds709
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.192 22.8795 11.238 23.0795 ;
 END
 END vccd_1p0.gds709
 PIN vccd_1p0.gds710
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.52 22.8795 10.566 23.0795 ;
 END
 END vccd_1p0.gds710
 PIN vccd_1p0.gds711
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.894 25.238 19.934 25.438 ;
 END
 END vccd_1p0.gds711
 PIN vccd_1p0.gds712
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.222 25.238 19.262 25.438 ;
 END
 END vccd_1p0.gds712
 PIN vccd_1p0.gds713
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.55 25.238 18.59 25.438 ;
 END
 END vccd_1p0.gds713
 PIN vccd_1p0.gds714
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.958 21.826 19.998 22.026 ;
 END
 END vccd_1p0.gds714
 PIN vccd_1p0.gds715
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.018 22.3645 17.074 22.5645 ;
 END
 END vccd_1p0.gds715
 PIN vccd_1p0.gds716
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.76 22.8795 19.806 23.0795 ;
 END
 END vccd_1p0.gds716
 PIN vccd_1p0.gds717
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.606 22.767 15.662 22.967 ;
 END
 END vccd_1p0.gds717
 PIN vccd_1p0.gds718
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 20.9415 15.742 21.1415 ;
 END
 END vccd_1p0.gds718
 PIN vccd_1p0.gds719
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 20.712 15.29 20.912 ;
 END
 END vccd_1p0.gds719
 PIN vccd_1p0.gds720
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 20.728 16.226 20.928 ;
 END
 END vccd_1p0.gds720
 PIN vccd_1p0.gds721
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 20.9905 17.574 21.1905 ;
 END
 END vccd_1p0.gds721
 PIN vccd_1p0.gds722
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 21.0135 17.154 21.2135 ;
 END
 END vccd_1p0.gds722
 PIN vccd_1p0.gds723
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 21.523 17.734 21.723 ;
 END
 END vccd_1p0.gds723
 PIN vccd_1p0.gds724
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 20.7045 15.498 20.9045 ;
 END
 END vccd_1p0.gds724
 PIN vccd_1p0.gds725
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.438 23.3685 17.494 23.5685 ;
 END
 END vccd_1p0.gds725
 PIN vccd_1p0.gds726
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.25 23.4885 16.31 23.6885 ;
 END
 END vccd_1p0.gds726
 PIN vccd_1p0.gds727
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.416 22.901 18.462 23.101 ;
 END
 END vccd_1p0.gds727
 PIN vccd_1p0.gds728
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.088 22.8795 19.134 23.0795 ;
 END
 END vccd_1p0.gds728
 PIN vccd_1p0.gds729
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.286 21.826 19.326 22.026 ;
 END
 END vccd_1p0.gds729
 PIN vccd_1p0.gds730
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.614 22.112 18.654 22.312 ;
 END
 END vccd_1p0.gds730
 PIN vccd_1p0.gds731
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.514 24.901 16.57 25.101 ;
 END
 END vccd_1p0.gds731
 PIN vccd_1p0.gds732
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 22.962 17.962 23.162 ;
 END
 END vccd_1p0.gds732
 PIN vccd_1p0.gds733
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 22.6615 18.09 22.8615 ;
 END
 END vccd_1p0.gds733
 PIN vccd_1p0.gds734
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.018 25.238 25.058 25.438 ;
 END
 END vccd_1p0.gds734
 PIN vccd_1p0.gds735
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.346 25.362 24.386 25.562 ;
 END
 END vccd_1p0.gds735
 PIN vccd_1p0.gds736
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.254 25.238 23.294 25.438 ;
 END
 END vccd_1p0.gds736
 PIN vccd_1p0.gds737
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.582 25.238 22.622 25.438 ;
 END
 END vccd_1p0.gds737
 PIN vccd_1p0.gds738
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.91 25.238 21.95 25.438 ;
 END
 END vccd_1p0.gds738
 PIN vccd_1p0.gds739
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.238 25.238 21.278 25.438 ;
 END
 END vccd_1p0.gds739
 PIN vccd_1p0.gds740
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.566 25.238 20.606 25.438 ;
 END
 END vccd_1p0.gds740
 PIN vccd_1p0.gds741
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.082 21.826 25.122 22.026 ;
 END
 END vccd_1p0.gds741
 PIN vccd_1p0.gds742
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.41 21.8735 24.45 22.0735 ;
 END
 END vccd_1p0.gds742
 PIN vccd_1p0.gds743
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.318 22.112 23.358 22.312 ;
 END
 END vccd_1p0.gds743
 PIN vccd_1p0.gds744
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.646 21.826 22.686 22.026 ;
 END
 END vccd_1p0.gds744
 PIN vccd_1p0.gds745
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.974 21.826 22.014 22.026 ;
 END
 END vccd_1p0.gds745
 PIN vccd_1p0.gds746
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.302 21.826 21.342 22.026 ;
 END
 END vccd_1p0.gds746
 PIN vccd_1p0.gds747
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.63 21.826 20.67 22.026 ;
 END
 END vccd_1p0.gds747
 PIN vccd_1p0.gds748
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.884 22.8795 24.93 23.0795 ;
 END
 END vccd_1p0.gds748
 PIN vccd_1p0.gds749
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.212 22.901 24.258 23.101 ;
 END
 END vccd_1p0.gds749
 PIN vccd_1p0.gds750
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.12 22.968 23.166 23.168 ;
 END
 END vccd_1p0.gds750
 PIN vccd_1p0.gds751
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.448 22.8795 22.494 23.0795 ;
 END
 END vccd_1p0.gds751
 PIN vccd_1p0.gds752
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.776 22.8795 21.822 23.0795 ;
 END
 END vccd_1p0.gds752
 PIN vccd_1p0.gds753
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.104 22.8795 21.15 23.0795 ;
 END
 END vccd_1p0.gds753
 PIN vccd_1p0.gds754
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.432 22.8795 20.478 23.0795 ;
 END
 END vccd_1p0.gds754
 PIN vccd_1p0.gds755
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 22.7385 23.842 22.9385 ;
 END
 END vccd_1p0.gds755
 PIN vccd_1p0.gds756
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.05 25.238 29.09 25.438 ;
 END
 END vccd_1p0.gds756
 PIN vccd_1p0.gds757
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.378 25.238 28.418 25.438 ;
 END
 END vccd_1p0.gds757
 PIN vccd_1p0.gds758
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.706 25.238 27.746 25.438 ;
 END
 END vccd_1p0.gds758
 PIN vccd_1p0.gds759
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.034 25.238 27.074 25.438 ;
 END
 END vccd_1p0.gds759
 PIN vccd_1p0.gds760
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.362 25.238 26.402 25.438 ;
 END
 END vccd_1p0.gds760
 PIN vccd_1p0.gds761
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.69 25.238 25.73 25.438 ;
 END
 END vccd_1p0.gds761
 PIN vccd_1p0.gds762
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.114 21.8735 29.154 22.0735 ;
 END
 END vccd_1p0.gds762
 PIN vccd_1p0.gds763
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.442 21.826 28.482 22.026 ;
 END
 END vccd_1p0.gds763
 PIN vccd_1p0.gds764
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.77 21.826 27.81 22.026 ;
 END
 END vccd_1p0.gds764
 PIN vccd_1p0.gds765
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.098 21.826 27.138 22.026 ;
 END
 END vccd_1p0.gds765
 PIN vccd_1p0.gds766
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.426 21.826 26.466 22.026 ;
 END
 END vccd_1p0.gds766
 PIN vccd_1p0.gds767
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.754 21.826 25.794 22.026 ;
 END
 END vccd_1p0.gds767
 PIN vccd_1p0.gds768
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 24.432 30.19 24.632 ;
 END
 END vccd_1p0.gds768
 PIN vccd_1p0.gds769
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 24.056 29.706 24.256 ;
 END
 END vccd_1p0.gds769
 PIN vccd_1p0.gds770
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.916 22.8795 28.962 23.0795 ;
 END
 END vccd_1p0.gds770
 PIN vccd_1p0.gds771
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.244 22.8795 28.29 23.0795 ;
 END
 END vccd_1p0.gds771
 PIN vccd_1p0.gds772
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.572 22.8795 27.618 23.0795 ;
 END
 END vccd_1p0.gds772
 PIN vccd_1p0.gds773
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.9 22.8795 26.946 23.0795 ;
 END
 END vccd_1p0.gds773
 PIN vccd_1p0.gds774
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.228 22.8795 26.274 23.0795 ;
 END
 END vccd_1p0.gds774
 PIN vccd_1p0.gds775
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.556 22.8795 25.602 23.0795 ;
 END
 END vccd_1p0.gds775
 PIN vccd_1p0.gds776
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.73 22.434 29.77 22.634 ;
 END
 END vccd_1p0.gds776
 PIN vccd_1p0.gds777
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 20.984 29.95 21.184 ;
 END
 END vccd_1p0.gds777
 PIN vccd_1p0.gds778
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 20.737 29.578 20.937 ;
 END
 END vccd_1p0.gds778
 PIN vccd_1p0.gds779
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 23.3505 32.342 23.5505 ;
 END
 END vccd_1p0.gds779
 PIN vccd_1p0.gds780
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 22.7035 31.986 22.9035 ;
 END
 END vccd_1p0.gds780
 PIN vccd_1p0.gds781
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.314 21.013 30.37 21.213 ;
 END
 END vccd_1p0.gds781
 PIN vccd_1p0.gds782
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 21.573 31.03 21.773 ;
 END
 END vccd_1p0.gds782
 PIN vccd_1p0.gds783
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.658 22.767 32.714 22.967 ;
 END
 END vccd_1p0.gds783
 PIN vccd_1p0.gds784
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.302 23.4885 33.362 23.6885 ;
 END
 END vccd_1p0.gds784
 PIN vccd_1p0.gds785
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.49 23.3685 34.546 23.5685 ;
 END
 END vccd_1p0.gds785
 PIN vccd_1p0.gds786
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.566 24.901 33.622 25.101 ;
 END
 END vccd_1p0.gds786
 PIN vccd_1p0.gds787
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 20.728 33.278 20.928 ;
 END
 END vccd_1p0.gds787
 PIN vccd_1p0.gds788
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 20.738 30.79 20.938 ;
 END
 END vccd_1p0.gds788
 PIN vccd_1p0.gds789
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 20.712 32.342 20.912 ;
 END
 END vccd_1p0.gds789
 PIN vccd_1p0.gds790
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 20.5055 31.986 20.7055 ;
 END
 END vccd_1p0.gds790
 PIN vccd_1p0.gds791
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 20.9785 31.794 21.1785 ;
 END
 END vccd_1p0.gds791
 PIN vccd_1p0.gds792
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 20.9905 34.626 21.1905 ;
 END
 END vccd_1p0.gds792
 PIN vccd_1p0.gds793
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 22.6615 35.142 22.8615 ;
 END
 END vccd_1p0.gds793
 PIN vccd_1p0.gds794
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 22.962 35.014 23.162 ;
 END
 END vccd_1p0.gds794
 PIN vccd_1p0.gds795
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 21.0135 34.206 21.2135 ;
 END
 END vccd_1p0.gds795
 PIN vccd_1p0.gds796
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 20.9415 32.794 21.1415 ;
 END
 END vccd_1p0.gds796
 PIN vccd_1p0.gds797
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 20.7045 32.55 20.9045 ;
 END
 END vccd_1p0.gds797
 PIN vccd_1p0.gds798
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 21.523 34.786 21.723 ;
 END
 END vccd_1p0.gds798
 PIN vccd_1p0.gds799
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.07 22.3645 34.126 22.5645 ;
 END
 END vccd_1p0.gds799
 PIN vccd_1p0.gds800
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.634 25.238 39.674 25.438 ;
 END
 END vccd_1p0.gds800
 PIN vccd_1p0.gds801
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.962 25.238 39.002 25.438 ;
 END
 END vccd_1p0.gds801
 PIN vccd_1p0.gds802
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.29 25.238 38.33 25.438 ;
 END
 END vccd_1p0.gds802
 PIN vccd_1p0.gds803
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.618 25.238 37.658 25.438 ;
 END
 END vccd_1p0.gds803
 PIN vccd_1p0.gds804
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.946 25.238 36.986 25.438 ;
 END
 END vccd_1p0.gds804
 PIN vccd_1p0.gds805
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.274 25.238 36.314 25.438 ;
 END
 END vccd_1p0.gds805
 PIN vccd_1p0.gds806
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.602 25.238 35.642 25.438 ;
 END
 END vccd_1p0.gds806
 PIN vccd_1p0.gds807
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.468 22.901 35.514 23.101 ;
 END
 END vccd_1p0.gds807
 PIN vccd_1p0.gds808
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.172 22.968 40.218 23.168 ;
 END
 END vccd_1p0.gds808
 PIN vccd_1p0.gds809
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.5 22.8795 39.546 23.0795 ;
 END
 END vccd_1p0.gds809
 PIN vccd_1p0.gds810
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.698 21.826 39.738 22.026 ;
 END
 END vccd_1p0.gds810
 PIN vccd_1p0.gds811
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.828 22.8795 38.874 23.0795 ;
 END
 END vccd_1p0.gds811
 PIN vccd_1p0.gds812
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.026 21.826 39.066 22.026 ;
 END
 END vccd_1p0.gds812
 PIN vccd_1p0.gds813
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.156 22.8795 38.202 23.0795 ;
 END
 END vccd_1p0.gds813
 PIN vccd_1p0.gds814
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.354 21.826 38.394 22.026 ;
 END
 END vccd_1p0.gds814
 PIN vccd_1p0.gds815
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.484 22.8795 37.53 23.0795 ;
 END
 END vccd_1p0.gds815
 PIN vccd_1p0.gds816
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.682 21.826 37.722 22.026 ;
 END
 END vccd_1p0.gds816
 PIN vccd_1p0.gds817
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.812 22.8795 36.858 23.0795 ;
 END
 END vccd_1p0.gds817
 PIN vccd_1p0.gds818
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.01 21.826 37.05 22.026 ;
 END
 END vccd_1p0.gds818
 PIN vccd_1p0.gds819
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.14 22.8795 36.186 23.0795 ;
 END
 END vccd_1p0.gds819
 PIN vccd_1p0.gds820
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.338 21.826 36.378 22.026 ;
 END
 END vccd_1p0.gds820
 PIN vccd_1p0.gds821
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.666 22.112 35.706 22.312 ;
 END
 END vccd_1p0.gds821
 PIN vccd_1p0.gds822
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.758 25.238 44.798 25.438 ;
 END
 END vccd_1p0.gds822
 PIN vccd_1p0.gds823
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.086 25.238 44.126 25.438 ;
 END
 END vccd_1p0.gds823
 PIN vccd_1p0.gds824
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.414 25.238 43.454 25.438 ;
 END
 END vccd_1p0.gds824
 PIN vccd_1p0.gds825
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.742 25.238 42.782 25.438 ;
 END
 END vccd_1p0.gds825
 PIN vccd_1p0.gds826
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.07 25.238 42.11 25.438 ;
 END
 END vccd_1p0.gds826
 PIN vccd_1p0.gds827
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.398 25.362 41.438 25.562 ;
 END
 END vccd_1p0.gds827
 PIN vccd_1p0.gds828
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.306 25.238 40.346 25.438 ;
 END
 END vccd_1p0.gds828
 PIN vccd_1p0.gds829
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.296 22.8795 45.342 23.0795 ;
 END
 END vccd_1p0.gds829
 PIN vccd_1p0.gds830
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.624 22.8795 44.67 23.0795 ;
 END
 END vccd_1p0.gds830
 PIN vccd_1p0.gds831
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.822 21.826 44.862 22.026 ;
 END
 END vccd_1p0.gds831
 PIN vccd_1p0.gds832
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.952 22.8795 43.998 23.0795 ;
 END
 END vccd_1p0.gds832
 PIN vccd_1p0.gds833
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.15 21.826 44.19 22.026 ;
 END
 END vccd_1p0.gds833
 PIN vccd_1p0.gds834
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.28 22.8795 43.326 23.0795 ;
 END
 END vccd_1p0.gds834
 PIN vccd_1p0.gds835
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.478 21.826 43.518 22.026 ;
 END
 END vccd_1p0.gds835
 PIN vccd_1p0.gds836
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.608 22.8795 42.654 23.0795 ;
 END
 END vccd_1p0.gds836
 PIN vccd_1p0.gds837
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.806 21.826 42.846 22.026 ;
 END
 END vccd_1p0.gds837
 PIN vccd_1p0.gds838
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.936 22.8795 41.982 23.0795 ;
 END
 END vccd_1p0.gds838
 PIN vccd_1p0.gds839
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.134 21.826 42.174 22.026 ;
 END
 END vccd_1p0.gds839
 PIN vccd_1p0.gds840
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.264 22.901 41.31 23.101 ;
 END
 END vccd_1p0.gds840
 PIN vccd_1p0.gds841
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.462 21.8735 41.502 22.0735 ;
 END
 END vccd_1p0.gds841
 PIN vccd_1p0.gds842
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.37 22.112 40.41 22.312 ;
 END
 END vccd_1p0.gds842
 PIN vccd_1p0.gds843
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 22.7385 40.894 22.9385 ;
 END
 END vccd_1p0.gds843
 PIN vccd_1p0.gds844
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.102 25.238 46.142 25.438 ;
 END
 END vccd_1p0.gds844
 PIN vccd_1p0.gds845
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.43 25.238 45.47 25.438 ;
 END
 END vccd_1p0.gds845
 PIN vccd_1p0.gds846
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 24.432 47.242 24.632 ;
 END
 END vccd_1p0.gds846
 PIN vccd_1p0.gds847
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 24.056 46.758 24.256 ;
 END
 END vccd_1p0.gds847
 PIN vccd_1p0.gds848
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 23.3505 49.394 23.5505 ;
 END
 END vccd_1p0.gds848
 PIN vccd_1p0.gds849
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 22.7035 49.038 22.9035 ;
 END
 END vccd_1p0.gds849
 PIN vccd_1p0.gds850
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.782 22.434 46.822 22.634 ;
 END
 END vccd_1p0.gds850
 PIN vccd_1p0.gds851
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.968 22.8795 46.014 23.0795 ;
 END
 END vccd_1p0.gds851
 PIN vccd_1p0.gds852
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.166 21.8735 46.206 22.0735 ;
 END
 END vccd_1p0.gds852
 PIN vccd_1p0.gds853
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.494 21.826 45.534 22.026 ;
 END
 END vccd_1p0.gds853
 PIN vccd_1p0.gds854
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.366 21.013 47.422 21.213 ;
 END
 END vccd_1p0.gds854
 PIN vccd_1p0.gds855
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 21.573 48.082 21.773 ;
 END
 END vccd_1p0.gds855
 PIN vccd_1p0.gds856
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.71 22.767 49.766 22.967 ;
 END
 END vccd_1p0.gds856
 PIN vccd_1p0.gds857
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 20.738 47.842 20.938 ;
 END
 END vccd_1p0.gds857
 PIN vccd_1p0.gds858
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 20.712 49.394 20.912 ;
 END
 END vccd_1p0.gds858
 PIN vccd_1p0.gds859
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 20.5055 49.038 20.7055 ;
 END
 END vccd_1p0.gds859
 PIN vccd_1p0.gds860
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 20.9785 48.846 21.1785 ;
 END
 END vccd_1p0.gds860
 PIN vccd_1p0.gds861
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 20.9415 49.846 21.1415 ;
 END
 END vccd_1p0.gds861
 PIN vccd_1p0.gds862
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 20.7045 49.602 20.9045 ;
 END
 END vccd_1p0.gds862
 PIN vccd_1p0.gds863
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 20.984 47.002 21.184 ;
 END
 END vccd_1p0.gds863
 PIN vccd_1p0.gds864
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 20.737 46.63 20.937 ;
 END
 END vccd_1p0.gds864
 PIN vccd_1p0.gds865
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.67 25.238 54.71 25.438 ;
 END
 END vccd_1p0.gds865
 PIN vccd_1p0.gds866
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.998 25.238 54.038 25.438 ;
 END
 END vccd_1p0.gds866
 PIN vccd_1p0.gds867
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.326 25.238 53.366 25.438 ;
 END
 END vccd_1p0.gds867
 PIN vccd_1p0.gds868
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.654 25.238 52.694 25.438 ;
 END
 END vccd_1p0.gds868
 PIN vccd_1p0.gds869
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.354 23.4885 50.414 23.6885 ;
 END
 END vccd_1p0.gds869
 PIN vccd_1p0.gds870
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.542 23.3685 51.598 23.5685 ;
 END
 END vccd_1p0.gds870
 PIN vccd_1p0.gds871
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.618 24.901 50.674 25.101 ;
 END
 END vccd_1p0.gds871
 PIN vccd_1p0.gds872
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.52 22.901 52.566 23.101 ;
 END
 END vccd_1p0.gds872
 PIN vccd_1p0.gds873
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.208 22.8795 55.254 23.0795 ;
 END
 END vccd_1p0.gds873
 PIN vccd_1p0.gds874
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.536 22.8795 54.582 23.0795 ;
 END
 END vccd_1p0.gds874
 PIN vccd_1p0.gds875
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.734 21.826 54.774 22.026 ;
 END
 END vccd_1p0.gds875
 PIN vccd_1p0.gds876
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.864 22.8795 53.91 23.0795 ;
 END
 END vccd_1p0.gds876
 PIN vccd_1p0.gds877
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.062 21.826 54.102 22.026 ;
 END
 END vccd_1p0.gds877
 PIN vccd_1p0.gds878
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 20.728 50.33 20.928 ;
 END
 END vccd_1p0.gds878
 PIN vccd_1p0.gds879
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 20.9905 51.678 21.1905 ;
 END
 END vccd_1p0.gds879
 PIN vccd_1p0.gds880
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 22.6615 52.194 22.8615 ;
 END
 END vccd_1p0.gds880
 PIN vccd_1p0.gds881
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 22.962 52.066 23.162 ;
 END
 END vccd_1p0.gds881
 PIN vccd_1p0.gds882
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 21.0135 51.258 21.2135 ;
 END
 END vccd_1p0.gds882
 PIN vccd_1p0.gds883
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 21.523 51.838 21.723 ;
 END
 END vccd_1p0.gds883
 PIN vccd_1p0.gds884
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.122 22.3645 51.178 22.5645 ;
 END
 END vccd_1p0.gds884
 PIN vccd_1p0.gds885
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.192 22.8795 53.238 23.0795 ;
 END
 END vccd_1p0.gds885
 PIN vccd_1p0.gds886
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.39 21.826 53.43 22.026 ;
 END
 END vccd_1p0.gds886
 PIN vccd_1p0.gds887
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.718 22.112 52.758 22.312 ;
 END
 END vccd_1p0.gds887
 PIN vccd_1p0.gds888
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.794 25.238 59.834 25.438 ;
 END
 END vccd_1p0.gds888
 PIN vccd_1p0.gds889
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.122 25.238 59.162 25.438 ;
 END
 END vccd_1p0.gds889
 PIN vccd_1p0.gds890
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.686 25.238 56.726 25.438 ;
 END
 END vccd_1p0.gds890
 PIN vccd_1p0.gds891
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.014 25.238 56.054 25.438 ;
 END
 END vccd_1p0.gds891
 PIN vccd_1p0.gds892
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.342 25.238 55.382 25.438 ;
 END
 END vccd_1p0.gds892
 PIN vccd_1p0.gds893
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.45 25.362 58.49 25.562 ;
 END
 END vccd_1p0.gds893
 PIN vccd_1p0.gds894
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.358 25.238 57.398 25.438 ;
 END
 END vccd_1p0.gds894
 PIN vccd_1p0.gds895
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.66 22.8795 59.706 23.0795 ;
 END
 END vccd_1p0.gds895
 PIN vccd_1p0.gds896
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.858 21.826 59.898 22.026 ;
 END
 END vccd_1p0.gds896
 PIN vccd_1p0.gds897
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.988 22.8795 59.034 23.0795 ;
 END
 END vccd_1p0.gds897
 PIN vccd_1p0.gds898
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.186 21.826 59.226 22.026 ;
 END
 END vccd_1p0.gds898
 PIN vccd_1p0.gds899
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.316 22.901 58.362 23.101 ;
 END
 END vccd_1p0.gds899
 PIN vccd_1p0.gds900
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.514 21.8735 58.554 22.0735 ;
 END
 END vccd_1p0.gds900
 PIN vccd_1p0.gds901
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.224 22.968 57.27 23.168 ;
 END
 END vccd_1p0.gds901
 PIN vccd_1p0.gds902
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.422 22.112 57.462 22.312 ;
 END
 END vccd_1p0.gds902
 PIN vccd_1p0.gds903
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.552 22.8795 56.598 23.0795 ;
 END
 END vccd_1p0.gds903
 PIN vccd_1p0.gds904
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.75 21.826 56.79 22.026 ;
 END
 END vccd_1p0.gds904
 PIN vccd_1p0.gds905
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.88 22.8795 55.926 23.0795 ;
 END
 END vccd_1p0.gds905
 PIN vccd_1p0.gds906
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.078 21.826 56.118 22.026 ;
 END
 END vccd_1p0.gds906
 PIN vccd_1p0.gds907
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.406 21.826 55.446 22.026 ;
 END
 END vccd_1p0.gds907
 PIN vccd_1p0.gds908
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 22.7385 57.946 22.9385 ;
 END
 END vccd_1p0.gds908
 PIN vccd_1p0.gds909
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.154 25.238 63.194 25.438 ;
 END
 END vccd_1p0.gds909
 PIN vccd_1p0.gds910
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.482 25.238 62.522 25.438 ;
 END
 END vccd_1p0.gds910
 PIN vccd_1p0.gds911
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.81 25.238 61.85 25.438 ;
 END
 END vccd_1p0.gds911
 PIN vccd_1p0.gds912
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.138 25.238 61.178 25.438 ;
 END
 END vccd_1p0.gds912
 PIN vccd_1p0.gds913
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.466 25.238 60.506 25.438 ;
 END
 END vccd_1p0.gds913
 PIN vccd_1p0.gds914
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 24.432 64.294 24.632 ;
 END
 END vccd_1p0.gds914
 PIN vccd_1p0.gds915
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 24.056 63.81 24.256 ;
 END
 END vccd_1p0.gds915
 PIN vccd_1p0.gds916
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.834 22.434 63.874 22.634 ;
 END
 END vccd_1p0.gds916
 PIN vccd_1p0.gds917
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.02 22.8795 63.066 23.0795 ;
 END
 END vccd_1p0.gds917
 PIN vccd_1p0.gds918
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.218 21.8735 63.258 22.0735 ;
 END
 END vccd_1p0.gds918
 PIN vccd_1p0.gds919
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.348 22.8795 62.394 23.0795 ;
 END
 END vccd_1p0.gds919
 PIN vccd_1p0.gds920
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.546 21.826 62.586 22.026 ;
 END
 END vccd_1p0.gds920
 PIN vccd_1p0.gds921
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.676 22.8795 61.722 23.0795 ;
 END
 END vccd_1p0.gds921
 PIN vccd_1p0.gds922
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.874 21.826 61.914 22.026 ;
 END
 END vccd_1p0.gds922
 PIN vccd_1p0.gds923
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.004 22.8795 61.05 23.0795 ;
 END
 END vccd_1p0.gds923
 PIN vccd_1p0.gds924
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.202 21.826 61.242 22.026 ;
 END
 END vccd_1p0.gds924
 PIN vccd_1p0.gds925
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.332 22.8795 60.378 23.0795 ;
 END
 END vccd_1p0.gds925
 PIN vccd_1p0.gds926
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.53 21.826 60.57 22.026 ;
 END
 END vccd_1p0.gds926
 PIN vccd_1p0.gds927
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.418 21.013 64.474 21.213 ;
 END
 END vccd_1p0.gds927
 PIN vccd_1p0.gds928
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 21.573 65.134 21.773 ;
 END
 END vccd_1p0.gds928
 PIN vccd_1p0.gds929
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 20.738 64.894 20.938 ;
 END
 END vccd_1p0.gds929
 PIN vccd_1p0.gds930
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 20.984 64.054 21.184 ;
 END
 END vccd_1p0.gds930
 PIN vccd_1p0.gds931
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 20.737 63.682 20.937 ;
 END
 END vccd_1p0.gds931
 PIN vccd_1p0.gds932
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.706 25.238 69.746 25.438 ;
 END
 END vccd_1p0.gds932
 PIN vccd_1p0.gds933
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 23.3505 66.446 23.5505 ;
 END
 END vccd_1p0.gds933
 PIN vccd_1p0.gds934
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 22.7035 66.09 22.9035 ;
 END
 END vccd_1p0.gds934
 PIN vccd_1p0.gds935
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.762 22.767 66.818 22.967 ;
 END
 END vccd_1p0.gds935
 PIN vccd_1p0.gds936
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.406 23.4885 67.466 23.6885 ;
 END
 END vccd_1p0.gds936
 PIN vccd_1p0.gds937
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.572 22.901 69.618 23.101 ;
 END
 END vccd_1p0.gds937
 PIN vccd_1p0.gds938
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 20.728 67.382 20.928 ;
 END
 END vccd_1p0.gds938
 PIN vccd_1p0.gds939
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 20.712 66.446 20.912 ;
 END
 END vccd_1p0.gds939
 PIN vccd_1p0.gds940
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 20.5055 66.09 20.7055 ;
 END
 END vccd_1p0.gds940
 PIN vccd_1p0.gds941
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 20.9785 65.898 21.1785 ;
 END
 END vccd_1p0.gds941
 PIN vccd_1p0.gds942
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 20.9905 68.73 21.1905 ;
 END
 END vccd_1p0.gds942
 PIN vccd_1p0.gds943
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 22.6615 69.246 22.8615 ;
 END
 END vccd_1p0.gds943
 PIN vccd_1p0.gds944
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 22.962 69.118 23.162 ;
 END
 END vccd_1p0.gds944
 PIN vccd_1p0.gds945
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 21.0135 68.31 21.2135 ;
 END
 END vccd_1p0.gds945
 PIN vccd_1p0.gds946
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 20.9415 66.898 21.1415 ;
 END
 END vccd_1p0.gds946
 PIN vccd_1p0.gds947
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 20.7045 66.654 20.9045 ;
 END
 END vccd_1p0.gds947
 PIN vccd_1p0.gds948
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 21.523 68.89 21.723 ;
 END
 END vccd_1p0.gds948
 PIN vccd_1p0.gds949
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.174 22.3645 68.23 22.5645 ;
 END
 END vccd_1p0.gds949
 PIN vccd_1p0.gds950
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.244 22.8795 70.29 23.0795 ;
 END
 END vccd_1p0.gds950
 PIN vccd_1p0.gds951
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.77 22.112 69.81 22.312 ;
 END
 END vccd_1p0.gds951
 PIN vccd_1p0.gds952
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.594 23.3685 68.65 23.5685 ;
 END
 END vccd_1p0.gds952
 PIN vccd_1p0.gds953
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.67 24.901 67.726 25.101 ;
 END
 END vccd_1p0.gds953
 PIN vccd_1p0.gds954
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.41 25.238 74.45 25.438 ;
 END
 END vccd_1p0.gds954
 PIN vccd_1p0.gds955
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.738 25.238 73.778 25.438 ;
 END
 END vccd_1p0.gds955
 PIN vccd_1p0.gds956
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.066 25.238 73.106 25.438 ;
 END
 END vccd_1p0.gds956
 PIN vccd_1p0.gds957
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.394 25.238 72.434 25.438 ;
 END
 END vccd_1p0.gds957
 PIN vccd_1p0.gds958
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.722 25.238 71.762 25.438 ;
 END
 END vccd_1p0.gds958
 PIN vccd_1p0.gds959
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.05 25.238 71.09 25.438 ;
 END
 END vccd_1p0.gds959
 PIN vccd_1p0.gds960
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.378 25.238 70.418 25.438 ;
 END
 END vccd_1p0.gds960
 PIN vccd_1p0.gds961
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.276 23.004 74.322 23.204 ;
 END
 END vccd_1p0.gds961
 PIN vccd_1p0.gds962
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.474 21.826 74.514 22.026 ;
 END
 END vccd_1p0.gds962
 PIN vccd_1p0.gds963
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.604 22.8795 73.65 23.0795 ;
 END
 END vccd_1p0.gds963
 PIN vccd_1p0.gds964
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.802 21.826 73.842 22.026 ;
 END
 END vccd_1p0.gds964
 PIN vccd_1p0.gds965
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.932 22.8795 72.978 23.0795 ;
 END
 END vccd_1p0.gds965
 PIN vccd_1p0.gds966
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.13 21.826 73.17 22.026 ;
 END
 END vccd_1p0.gds966
 PIN vccd_1p0.gds967
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.26 22.8795 72.306 23.0795 ;
 END
 END vccd_1p0.gds967
 PIN vccd_1p0.gds968
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.458 21.826 72.498 22.026 ;
 END
 END vccd_1p0.gds968
 PIN vccd_1p0.gds969
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.588 22.8795 71.634 23.0795 ;
 END
 END vccd_1p0.gds969
 PIN vccd_1p0.gds970
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.786 21.826 71.826 22.026 ;
 END
 END vccd_1p0.gds970
 PIN vccd_1p0.gds971
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.916 22.8795 70.962 23.0795 ;
 END
 END vccd_1p0.gds971
 PIN vccd_1p0.gds972
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.114 21.826 71.154 22.026 ;
 END
 END vccd_1p0.gds972
 PIN vccd_1p0.gds973
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.442 21.826 70.482 22.026 ;
 END
 END vccd_1p0.gds973
 PIN vccd_1p0.gds974
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 29.1795 0.43 29.3795 ;
 END
 END vccd_1p0.gds974
 PIN vccd_1p0.gds975
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 29.237 1.542 29.437 ;
 END
 END vccd_1p0.gds975
 PIN vccd_1p0.gds976
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 30.3795 5.202 30.5795 ;
 END
 END vccd_1p0.gds976
 PIN vccd_1p0.gds977
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 27.977 0.548 28.177 ;
 END
 END vccd_1p0.gds977
 PIN vccd_1p0.gds978
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 27.1995 1.542 27.3995 ;
 END
 END vccd_1p0.gds978
 PIN vccd_1p0.gds979
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 26.712 2.462 26.912 ;
 END
 END vccd_1p0.gds979
 PIN vccd_1p0.gds980
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 29.47 1.782 29.67 ;
 END
 END vccd_1p0.gds980
 PIN vccd_1p0.gds981
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 28.0455 0.858 28.2455 ;
 END
 END vccd_1p0.gds981
 PIN vccd_1p0.gds982
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 27.883 1.362 28.083 ;
 END
 END vccd_1p0.gds982
 PIN vccd_1p0.gds983
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 27.9615 1.218 28.1615 ;
 END
 END vccd_1p0.gds983
 PIN vccd_1p0.gds984
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 27.962 1.09 28.162 ;
 END
 END vccd_1p0.gds984
 PIN vccd_1p0.gds985
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 29.928 2.202 30.128 ;
 END
 END vccd_1p0.gds985
 PIN vccd_1p0.gds986
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 27.653 2.622 27.853 ;
 END
 END vccd_1p0.gds986
 PIN vccd_1p0.gds987
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 30.3965 2.462 30.5965 ;
 END
 END vccd_1p0.gds987
 PIN vccd_1p0.gds988
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 27.867 3.042 28.067 ;
 END
 END vccd_1p0.gds988
 PIN vccd_1p0.gds989
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 27.2095 1.962 27.4095 ;
 END
 END vccd_1p0.gds989
 PIN vccd_1p0.gds990
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 27.9505 2.882 28.1505 ;
 END
 END vccd_1p0.gds990
 PIN vccd_1p0.gds991
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 27.793 3.39 27.993 ;
 END
 END vccd_1p0.gds991
 PIN vccd_1p0.gds992
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 28.0165 3.262 28.2165 ;
 END
 END vccd_1p0.gds992
 PIN vccd_1p0.gds993
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 28.612 5.202 28.812 ;
 END
 END vccd_1p0.gds993
 PIN vccd_1p0.gds994
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 26.812 4.258 27.012 ;
 END
 END vccd_1p0.gds994
 PIN vccd_1p0.gds995
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 27.916 3.858 28.116 ;
 END
 END vccd_1p0.gds995
 PIN vccd_1p0.gds996
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 27.817 4.546 28.017 ;
 END
 END vccd_1p0.gds996
 PIN vccd_1p0.gds997
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 27.606 5.01 27.806 ;
 END
 END vccd_1p0.gds997
 PIN vccd_1p0.gds998
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 4.34 29.452 4.396 29.652 ;
 RECT 4.76 29.428 4.816 29.628 ;
 RECT 5.096 29.452 5.152 29.652 ;
 RECT 3.584 29.2635 3.64 29.4635 ;
 RECT 4.172 29.3495 4.228 29.5495 ;
 RECT 4.928 29.306 4.984 29.506 ;
 END
 END vccd_1p0.gds998
 PIN vccd_1p0.gds999
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.566 25.8165 9.606 26.0165 ;
 END
 END vccd_1p0.gds999
 PIN vccd_1p0.gds1000
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.894 25.8165 8.934 26.0165 ;
 END
 END vccd_1p0.gds1000
 PIN vccd_1p0.gds1001
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.222 25.8165 8.262 26.0165 ;
 END
 END vccd_1p0.gds1001
 PIN vccd_1p0.gds1002
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.55 25.8165 7.59 26.0165 ;
 END
 END vccd_1p0.gds1002
 PIN vccd_1p0.gds1003
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.798 27.6555 9.858 27.8555 ;
 END
 END vccd_1p0.gds1003
 PIN vccd_1p0.gds1004
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.134 27.624 10.194 27.824 ;
 END
 END vccd_1p0.gds1004
 PIN vccd_1p0.gds1005
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.126 27.6555 9.186 27.8555 ;
 END
 END vccd_1p0.gds1005
 PIN vccd_1p0.gds1006
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 9.462 27.624 9.522 27.824 ;
 END
 END vccd_1p0.gds1006
 PIN vccd_1p0.gds1007
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.454 27.6555 8.514 27.8555 ;
 END
 END vccd_1p0.gds1007
 PIN vccd_1p0.gds1008
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.79 27.624 8.85 27.824 ;
 END
 END vccd_1p0.gds1008
 PIN vccd_1p0.gds1009
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.782 27.6555 7.842 27.8555 ;
 END
 END vccd_1p0.gds1009
 PIN vccd_1p0.gds1010
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 8.118 27.624 8.178 27.824 ;
 END
 END vccd_1p0.gds1010
 PIN vccd_1p0.gds1011
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.11 27.6555 7.17 27.8555 ;
 END
 END vccd_1p0.gds1011
 PIN vccd_1p0.gds1012
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 7.446 27.624 7.506 27.824 ;
 END
 END vccd_1p0.gds1012
 PIN vccd_1p0.gds1013
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 27.9055 6.838 28.1055 ;
 END
 END vccd_1p0.gds1013
 PIN vccd_1p0.gds1014
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 27.9205 5.602 28.1205 ;
 END
 END vccd_1p0.gds1014
 PIN vccd_1p0.gds1015
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 30.403 6.05 30.603 ;
 END
 END vccd_1p0.gds1015
 PIN vccd_1p0.gds1016
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 26.087 5.41 26.287 ;
 END
 END vccd_1p0.gds1016
 PIN vccd_1p0.gds1017
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 29.6505 5.922 29.8505 ;
 END
 END vccd_1p0.gds1017
 PIN vccd_1p0.gds1018
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 28.8225 6.306 29.0225 ;
 END
 END vccd_1p0.gds1018
 PIN vccd_1p0.gds1019
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 27.829 6.582 28.029 ;
 END
 END vccd_1p0.gds1019
 PIN vccd_1p0.gds1020
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 9.968 28.1755 10.024 28.3755 ;
 RECT 9.8 28.1455 9.856 28.3455 ;
 RECT 9.296 28.1755 9.352 28.3755 ;
 RECT 9.128 28.1455 9.184 28.3455 ;
 RECT 9.632 28.044 9.688 28.244 ;
 RECT 8.624 28.1755 8.68 28.3755 ;
 RECT 8.456 28.1455 8.512 28.3455 ;
 RECT 8.96 28.044 9.016 28.244 ;
 RECT 7.952 28.1755 8.008 28.3755 ;
 RECT 7.784 28.1455 7.84 28.3455 ;
 RECT 8.288 28.044 8.344 28.244 ;
 RECT 6.944 28.044 7 28.244 ;
 RECT 7.28 28.1755 7.336 28.3755 ;
 RECT 7.112 28.1455 7.168 28.3455 ;
 RECT 7.616 28.044 7.672 28.244 ;
 RECT 5.6 29.3495 5.656 29.5495 ;
 RECT 5.264 29.3495 5.32 29.5495 ;
 RECT 5.432 29.2635 5.488 29.4635 ;
 RECT 5.936 29.2635 5.992 29.4635 ;
 RECT 5.768 29.2635 5.824 29.4635 ;
 RECT 6.44 29.278 6.496 29.478 ;
 RECT 6.272 29.2635 6.328 29.4635 ;
 RECT 6.104 29.452 6.16 29.652 ;
 END
 END vccd_1p0.gds1020
 PIN vccd_1p0.gds1021
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 29.584 13.978 29.784 ;
 END
 END vccd_1p0.gds1021
 PIN vccd_1p0.gds1022
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 27.777 14.398 27.977 ;
 END
 END vccd_1p0.gds1022
 PIN vccd_1p0.gds1023
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 29.584 14.398 29.784 ;
 END
 END vccd_1p0.gds1023
 PIN vccd_1p0.gds1024
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 26.687 14.934 26.887 ;
 END
 END vccd_1p0.gds1024
 PIN vccd_1p0.gds1025
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 28.6325 13.738 28.8325 ;
 END
 END vccd_1p0.gds1025
 PIN vccd_1p0.gds1026
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 29.075 13.138 29.275 ;
 END
 END vccd_1p0.gds1026
 PIN vccd_1p0.gds1027
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 27.4215 12.898 27.6215 ;
 END
 END vccd_1p0.gds1027
 PIN vccd_1p0.gds1028
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 28.1475 12.654 28.3475 ;
 END
 END vccd_1p0.gds1028
 PIN vccd_1p0.gds1029
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 26.8535 14.742 27.0535 ;
 END
 END vccd_1p0.gds1029
 PIN vccd_1p0.gds1030
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 28.351 13.978 28.551 ;
 END
 END vccd_1p0.gds1030
 PIN vccd_1p0.gds1031
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 25.533 13.978 25.733 ;
 END
 END vccd_1p0.gds1031
 PIN vccd_1p0.gds1032
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 29.7115 14.934 29.9115 ;
 END
 END vccd_1p0.gds1032
 PIN vccd_1p0.gds1033
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.254 25.8205 12.294 26.0205 ;
 END
 END vccd_1p0.gds1033
 PIN vccd_1p0.gds1034
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.582 25.8165 11.622 26.0165 ;
 END
 END vccd_1p0.gds1034
 PIN vccd_1p0.gds1035
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.91 25.8165 10.95 26.0165 ;
 END
 END vccd_1p0.gds1035
 PIN vccd_1p0.gds1036
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.238 25.8165 10.278 26.0165 ;
 END
 END vccd_1p0.gds1036
 PIN vccd_1p0.gds1037
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.814 27.6555 11.874 27.8555 ;
 END
 END vccd_1p0.gds1037
 PIN vccd_1p0.gds1038
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.15 27.624 12.21 27.824 ;
 END
 END vccd_1p0.gds1038
 PIN vccd_1p0.gds1039
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.142 27.6555 11.202 27.8555 ;
 END
 END vccd_1p0.gds1039
 PIN vccd_1p0.gds1040
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 11.478 27.624 11.538 27.824 ;
 END
 END vccd_1p0.gds1040
 PIN vccd_1p0.gds1041
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.47 27.6555 10.53 27.8555 ;
 END
 END vccd_1p0.gds1041
 PIN vccd_1p0.gds1042
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 10.806 27.624 10.866 27.824 ;
 END
 END vccd_1p0.gds1042
 PIN vccd_1p0.gds1043
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 12.74 27.6745 12.796 27.8745 ;
 RECT 13.244 27.486 13.3 27.686 ;
 RECT 12.572 27.76 12.628 27.96 ;
 RECT 15.092 27.76 15.148 27.96 ;
 RECT 14.924 27.854 14.98 28.054 ;
 RECT 14.756 27.6745 14.812 27.8745 ;
 RECT 14.588 27.6745 14.644 27.8745 ;
 RECT 14.42 27.6745 14.476 27.8745 ;
 RECT 14.252 27.6745 14.308 27.8745 ;
 RECT 14.084 27.76 14.14 27.96 ;
 RECT 13.916 27.854 13.972 28.054 ;
 RECT 13.748 27.6745 13.804 27.8745 ;
 RECT 11.984 28.1755 12.04 28.3755 ;
 RECT 11.816 28.1455 11.872 28.3455 ;
 RECT 12.32 28.044 12.376 28.244 ;
 RECT 11.312 28.1755 11.368 28.3755 ;
 RECT 11.144 28.1455 11.2 28.3455 ;
 RECT 11.648 28.044 11.704 28.244 ;
 RECT 10.64 28.1755 10.696 28.3755 ;
 RECT 10.472 28.1455 10.528 28.3455 ;
 RECT 10.976 28.044 11.032 28.244 ;
 RECT 10.304 28.044 10.36 28.244 ;
 END
 END vccd_1p0.gds1043
 PIN vccd_1p0.gds1044
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.71 27.6555 19.77 27.8555 ;
 END
 END vccd_1p0.gds1044
 PIN vccd_1p0.gds1045
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.046 27.624 20.106 27.824 ;
 END
 END vccd_1p0.gds1045
 PIN vccd_1p0.gds1046
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.334 27.875 16.39 28.075 ;
 END
 END vccd_1p0.gds1046
 PIN vccd_1p0.gds1047
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.15 25.8165 20.19 26.0165 ;
 END
 END vccd_1p0.gds1047
 PIN vccd_1p0.gds1048
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.478 25.8165 19.518 26.0165 ;
 END
 END vccd_1p0.gds1048
 PIN vccd_1p0.gds1049
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 29.648 16.226 29.848 ;
 END
 END vccd_1p0.gds1049
 PIN vccd_1p0.gds1050
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 28.28 15.742 28.48 ;
 END
 END vccd_1p0.gds1050
 PIN vccd_1p0.gds1051
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 29.516 15.29 29.716 ;
 END
 END vccd_1p0.gds1051
 PIN vccd_1p0.gds1052
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 25.982 17.962 26.182 ;
 END
 END vccd_1p0.gds1052
 PIN vccd_1p0.gds1053
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 27.5675 17.574 27.7675 ;
 END
 END vccd_1p0.gds1053
 PIN vccd_1p0.gds1054
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 29.679 18.09 29.879 ;
 END
 END vccd_1p0.gds1054
 PIN vccd_1p0.gds1055
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 29.5635 17.962 29.7635 ;
 END
 END vccd_1p0.gds1055
 PIN vccd_1p0.gds1056
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 29.4455 17.734 29.6455 ;
 END
 END vccd_1p0.gds1056
 PIN vccd_1p0.gds1057
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 28.0055 15.498 28.2055 ;
 END
 END vccd_1p0.gds1057
 PIN vccd_1p0.gds1058
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.806 25.8165 18.846 26.0165 ;
 END
 END vccd_1p0.gds1058
 PIN vccd_1p0.gds1059
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 25.9095 18.09 26.1095 ;
 END
 END vccd_1p0.gds1059
 PIN vccd_1p0.gds1060
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 27.2115 16.226 27.4115 ;
 END
 END vccd_1p0.gds1060
 PIN vccd_1p0.gds1061
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 27.223 17.154 27.423 ;
 END
 END vccd_1p0.gds1061
 PIN vccd_1p0.gds1062
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.038 27.6555 19.098 27.8555 ;
 END
 END vccd_1p0.gds1062
 PIN vccd_1p0.gds1063
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 19.374 27.624 19.434 27.824 ;
 END
 END vccd_1p0.gds1063
 PIN vccd_1p0.gds1064
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.366 27.5315 18.426 27.7315 ;
 END
 END vccd_1p0.gds1064
 PIN vccd_1p0.gds1065
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.702 27.624 18.762 27.824 ;
 END
 END vccd_1p0.gds1065
 PIN vccd_1p0.gds1066
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 19.88 28.1755 19.936 28.3755 ;
 RECT 19.712 28.1455 19.768 28.3455 ;
 RECT 20.216 28.044 20.272 28.244 ;
 RECT 15.26 27.76 15.316 27.96 ;
 RECT 15.428 27.76 15.484 27.96 ;
 RECT 17.276 27.76 17.332 27.96 ;
 RECT 17.108 27.76 17.164 27.96 ;
 RECT 15.596 27.6745 15.652 27.8745 ;
 RECT 17.612 27.6745 17.668 27.8745 ;
 RECT 17.444 27.6745 17.5 27.8745 ;
 RECT 17.948 27.5775 18.004 27.7775 ;
 RECT 19.208 28.1755 19.264 28.3755 ;
 RECT 19.04 28.1455 19.096 28.3455 ;
 RECT 19.544 28.044 19.6 28.244 ;
 RECT 18.536 28.1755 18.592 28.3755 ;
 RECT 18.2 28.044 18.256 28.244 ;
 RECT 18.368 28.1455 18.424 28.3455 ;
 RECT 18.872 28.044 18.928 28.244 ;
 RECT 17.78 27.76 17.836 27.96 ;
 END
 END vccd_1p0.gds1066
 PIN vccd_1p0.gds1067
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.834 27.6555 24.894 27.8555 ;
 END
 END vccd_1p0.gds1067
 PIN vccd_1p0.gds1068
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.17 27.624 25.23 27.824 ;
 END
 END vccd_1p0.gds1068
 PIN vccd_1p0.gds1069
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.162 27.6555 24.222 27.8555 ;
 END
 END vccd_1p0.gds1069
 PIN vccd_1p0.gds1070
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.498 27.624 24.558 27.824 ;
 END
 END vccd_1p0.gds1070
 PIN vccd_1p0.gds1071
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.07 27.6555 23.13 27.8555 ;
 END
 END vccd_1p0.gds1071
 PIN vccd_1p0.gds1072
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.406 27.624 23.466 27.824 ;
 END
 END vccd_1p0.gds1072
 PIN vccd_1p0.gds1073
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.398 27.6555 22.458 27.8555 ;
 END
 END vccd_1p0.gds1073
 PIN vccd_1p0.gds1074
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.734 27.624 22.794 27.824 ;
 END
 END vccd_1p0.gds1074
 PIN vccd_1p0.gds1075
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.726 27.6555 21.786 27.8555 ;
 END
 END vccd_1p0.gds1075
 PIN vccd_1p0.gds1076
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.062 27.624 22.122 27.824 ;
 END
 END vccd_1p0.gds1076
 PIN vccd_1p0.gds1077
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.054 27.6555 21.114 27.8555 ;
 END
 END vccd_1p0.gds1077
 PIN vccd_1p0.gds1078
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.39 27.624 21.45 27.824 ;
 END
 END vccd_1p0.gds1078
 PIN vccd_1p0.gds1079
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.382 27.6555 20.442 27.8555 ;
 END
 END vccd_1p0.gds1079
 PIN vccd_1p0.gds1080
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.718 27.624 20.778 27.824 ;
 END
 END vccd_1p0.gds1080
 PIN vccd_1p0.gds1081
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.838 25.8165 22.878 26.0165 ;
 END
 END vccd_1p0.gds1081
 PIN vccd_1p0.gds1082
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 22.166 25.8165 22.206 26.0165 ;
 END
 END vccd_1p0.gds1082
 PIN vccd_1p0.gds1083
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 21.494 25.8165 21.534 26.0165 ;
 END
 END vccd_1p0.gds1083
 PIN vccd_1p0.gds1084
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 20.822 25.8165 20.862 26.0165 ;
 END
 END vccd_1p0.gds1084
 PIN vccd_1p0.gds1085
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 24.602 25.8165 24.642 26.0165 ;
 END
 END vccd_1p0.gds1085
 PIN vccd_1p0.gds1086
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.51 25.858 23.55 26.058 ;
 END
 END vccd_1p0.gds1086
 PIN vccd_1p0.gds1087
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 27.9515 23.842 28.1515 ;
 END
 END vccd_1p0.gds1087
 PIN vccd_1p0.gds1088
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 25.004 28.1755 25.06 28.3755 ;
 RECT 24.836 28.1455 24.892 28.3455 ;
 RECT 24.332 28.1755 24.388 28.3755 ;
 RECT 23.996 28.044 24.052 28.244 ;
 RECT 24.164 28.1455 24.22 28.3455 ;
 RECT 24.668 28.044 24.724 28.244 ;
 RECT 23.24 28.1755 23.296 28.3755 ;
 RECT 23.072 28.1455 23.128 28.3455 ;
 RECT 23.576 28.044 23.632 28.244 ;
 RECT 22.568 28.1755 22.624 28.3755 ;
 RECT 22.4 28.1455 22.456 28.3455 ;
 RECT 22.904 28.044 22.96 28.244 ;
 RECT 21.896 28.1755 21.952 28.3755 ;
 RECT 21.728 28.1455 21.784 28.3455 ;
 RECT 22.232 28.044 22.288 28.244 ;
 RECT 21.224 28.1755 21.28 28.3755 ;
 RECT 21.056 28.1455 21.112 28.3455 ;
 RECT 21.56 28.044 21.616 28.244 ;
 RECT 20.552 28.1755 20.608 28.3755 ;
 RECT 20.888 28.044 20.944 28.244 ;
 RECT 20.384 28.1455 20.44 28.3455 ;
 RECT 23.828 27.6745 23.884 27.8745 ;
 END
 END vccd_1p0.gds1088
 PIN vccd_1p0.gds1089
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.866 27.6555 28.926 27.8555 ;
 END
 END vccd_1p0.gds1089
 PIN vccd_1p0.gds1090
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.202 27.624 29.262 27.824 ;
 END
 END vccd_1p0.gds1090
 PIN vccd_1p0.gds1091
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.194 27.6555 28.254 27.8555 ;
 END
 END vccd_1p0.gds1091
 PIN vccd_1p0.gds1092
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.53 27.624 28.59 27.824 ;
 END
 END vccd_1p0.gds1092
 PIN vccd_1p0.gds1093
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.522 27.6555 27.582 27.8555 ;
 END
 END vccd_1p0.gds1093
 PIN vccd_1p0.gds1094
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.858 27.624 27.918 27.824 ;
 END
 END vccd_1p0.gds1094
 PIN vccd_1p0.gds1095
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.85 27.6555 26.91 27.8555 ;
 END
 END vccd_1p0.gds1095
 PIN vccd_1p0.gds1096
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.186 27.624 27.246 27.824 ;
 END
 END vccd_1p0.gds1096
 PIN vccd_1p0.gds1097
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.178 27.6555 26.238 27.8555 ;
 END
 END vccd_1p0.gds1097
 PIN vccd_1p0.gds1098
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.514 27.624 26.574 27.824 ;
 END
 END vccd_1p0.gds1098
 PIN vccd_1p0.gds1099
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.506 27.6555 25.566 27.8555 ;
 END
 END vccd_1p0.gds1099
 PIN vccd_1p0.gds1100
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.842 27.624 25.902 27.824 ;
 END
 END vccd_1p0.gds1100
 PIN vccd_1p0.gds1101
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 28.634 25.8165 28.674 26.0165 ;
 END
 END vccd_1p0.gds1101
 PIN vccd_1p0.gds1102
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.962 25.8165 28.002 26.0165 ;
 END
 END vccd_1p0.gds1102
 PIN vccd_1p0.gds1103
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 27.29 25.8165 27.33 26.0165 ;
 END
 END vccd_1p0.gds1103
 PIN vccd_1p0.gds1104
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 26.618 25.8165 26.658 26.0165 ;
 END
 END vccd_1p0.gds1104
 PIN vccd_1p0.gds1105
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.946 25.8165 25.986 26.0165 ;
 END
 END vccd_1p0.gds1105
 PIN vccd_1p0.gds1106
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 25.274 25.8165 25.314 26.0165 ;
 END
 END vccd_1p0.gds1106
 PIN vccd_1p0.gds1107
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 28.1475 29.706 28.3475 ;
 END
 END vccd_1p0.gds1107
 PIN vccd_1p0.gds1108
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 27.4215 29.95 27.6215 ;
 END
 END vccd_1p0.gds1108
 PIN vccd_1p0.gds1109
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.306 25.8205 29.346 26.0205 ;
 END
 END vccd_1p0.gds1109
 PIN vccd_1p0.gds1110
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 29.036 28.1755 29.092 28.3755 ;
 RECT 28.868 28.1455 28.924 28.3455 ;
 RECT 29.372 28.044 29.428 28.244 ;
 RECT 28.364 28.1755 28.42 28.3755 ;
 RECT 28.196 28.1455 28.252 28.3455 ;
 RECT 28.7 28.044 28.756 28.244 ;
 RECT 27.692 28.1755 27.748 28.3755 ;
 RECT 27.524 28.1455 27.58 28.3455 ;
 RECT 28.028 28.044 28.084 28.244 ;
 RECT 27.02 28.1755 27.076 28.3755 ;
 RECT 26.852 28.1455 26.908 28.3455 ;
 RECT 27.356 28.044 27.412 28.244 ;
 RECT 26.348 28.1755 26.404 28.3755 ;
 RECT 26.18 28.1455 26.236 28.3455 ;
 RECT 26.684 28.044 26.74 28.244 ;
 RECT 25.676 28.1755 25.732 28.3755 ;
 RECT 25.508 28.1455 25.564 28.3455 ;
 RECT 26.012 28.044 26.068 28.244 ;
 RECT 25.34 28.044 25.396 28.244 ;
 RECT 29.792 27.6745 29.848 27.8745 ;
 RECT 29.624 27.76 29.68 27.96 ;
 END
 END vccd_1p0.gds1110
 PIN vccd_1p0.gds1111
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 29.584 31.03 29.784 ;
 END
 END vccd_1p0.gds1111
 PIN vccd_1p0.gds1112
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 27.777 31.45 27.977 ;
 END
 END vccd_1p0.gds1112
 PIN vccd_1p0.gds1113
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 29.648 33.278 29.848 ;
 END
 END vccd_1p0.gds1113
 PIN vccd_1p0.gds1114
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 29.584 31.45 29.784 ;
 END
 END vccd_1p0.gds1114
 PIN vccd_1p0.gds1115
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 25.9095 35.142 26.1095 ;
 END
 END vccd_1p0.gds1115
 PIN vccd_1p0.gds1116
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 25.982 35.014 26.182 ;
 END
 END vccd_1p0.gds1116
 PIN vccd_1p0.gds1117
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 29.516 32.342 29.716 ;
 END
 END vccd_1p0.gds1117
 PIN vccd_1p0.gds1118
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 28.6325 30.79 28.8325 ;
 END
 END vccd_1p0.gds1118
 PIN vccd_1p0.gds1119
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 29.075 30.19 29.275 ;
 END
 END vccd_1p0.gds1119
 PIN vccd_1p0.gds1120
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 25.533 31.03 25.733 ;
 END
 END vccd_1p0.gds1120
 PIN vccd_1p0.gds1121
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 28.351 31.03 28.551 ;
 END
 END vccd_1p0.gds1121
 PIN vccd_1p0.gds1122
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 26.687 31.986 26.887 ;
 END
 END vccd_1p0.gds1122
 PIN vccd_1p0.gds1123
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 26.8535 31.794 27.0535 ;
 END
 END vccd_1p0.gds1123
 PIN vccd_1p0.gds1124
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 27.5675 34.626 27.7675 ;
 END
 END vccd_1p0.gds1124
 PIN vccd_1p0.gds1125
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 29.679 35.142 29.879 ;
 END
 END vccd_1p0.gds1125
 PIN vccd_1p0.gds1126
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 29.5635 35.014 29.7635 ;
 END
 END vccd_1p0.gds1126
 PIN vccd_1p0.gds1127
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 27.223 34.206 27.423 ;
 END
 END vccd_1p0.gds1127
 PIN vccd_1p0.gds1128
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 28.0055 32.55 28.2055 ;
 END
 END vccd_1p0.gds1128
 PIN vccd_1p0.gds1129
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 29.7115 31.986 29.9115 ;
 END
 END vccd_1p0.gds1129
 PIN vccd_1p0.gds1130
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 29.4455 34.786 29.6455 ;
 END
 END vccd_1p0.gds1130
 PIN vccd_1p0.gds1131
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 28.28 32.794 28.48 ;
 END
 END vccd_1p0.gds1131
 PIN vccd_1p0.gds1132
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.386 27.875 33.442 28.075 ;
 END
 END vccd_1p0.gds1132
 PIN vccd_1p0.gds1133
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 27.2115 33.278 27.4115 ;
 END
 END vccd_1p0.gds1133
 PIN vccd_1p0.gds1134
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 32.312 27.76 32.368 27.96 ;
 RECT 30.296 27.486 30.352 27.686 ;
 RECT 32.144 27.76 32.2 27.96 ;
 RECT 31.976 27.854 32.032 28.054 ;
 RECT 31.808 27.6745 31.864 27.8745 ;
 RECT 31.64 27.6745 31.696 27.8745 ;
 RECT 31.472 27.6745 31.528 27.8745 ;
 RECT 31.304 27.6745 31.36 27.8745 ;
 RECT 31.136 27.76 31.192 27.96 ;
 RECT 30.968 27.854 31.024 28.054 ;
 RECT 30.8 27.6745 30.856 27.8745 ;
 RECT 32.648 27.6745 32.704 27.8745 ;
 RECT 32.48 27.76 32.536 27.96 ;
 RECT 35 27.5775 35.056 27.7775 ;
 RECT 34.832 27.76 34.888 27.96 ;
 RECT 34.664 27.6745 34.72 27.8745 ;
 RECT 34.496 27.6745 34.552 27.8745 ;
 RECT 34.328 27.76 34.384 27.96 ;
 RECT 34.16 27.76 34.216 27.96 ;
 END
 END vccd_1p0.gds1134
 PIN vccd_1p0.gds1135
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.122 27.6555 40.182 27.8555 ;
 END
 END vccd_1p0.gds1135
 PIN vccd_1p0.gds1136
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.45 27.6555 39.51 27.8555 ;
 END
 END vccd_1p0.gds1136
 PIN vccd_1p0.gds1137
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.786 27.624 39.846 27.824 ;
 END
 END vccd_1p0.gds1137
 PIN vccd_1p0.gds1138
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.778 27.6555 38.838 27.8555 ;
 END
 END vccd_1p0.gds1138
 PIN vccd_1p0.gds1139
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.114 27.624 39.174 27.824 ;
 END
 END vccd_1p0.gds1139
 PIN vccd_1p0.gds1140
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.106 27.6555 38.166 27.8555 ;
 END
 END vccd_1p0.gds1140
 PIN vccd_1p0.gds1141
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.442 27.624 38.502 27.824 ;
 END
 END vccd_1p0.gds1141
 PIN vccd_1p0.gds1142
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.434 27.6555 37.494 27.8555 ;
 END
 END vccd_1p0.gds1142
 PIN vccd_1p0.gds1143
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.77 27.624 37.83 27.824 ;
 END
 END vccd_1p0.gds1143
 PIN vccd_1p0.gds1144
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.762 27.6555 36.822 27.8555 ;
 END
 END vccd_1p0.gds1144
 PIN vccd_1p0.gds1145
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.098 27.624 37.158 27.824 ;
 END
 END vccd_1p0.gds1145
 PIN vccd_1p0.gds1146
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.09 27.6555 36.15 27.8555 ;
 END
 END vccd_1p0.gds1146
 PIN vccd_1p0.gds1147
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.426 27.624 36.486 27.824 ;
 END
 END vccd_1p0.gds1147
 PIN vccd_1p0.gds1148
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.418 27.5315 35.478 27.7315 ;
 END
 END vccd_1p0.gds1148
 PIN vccd_1p0.gds1149
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.754 27.624 35.814 27.824 ;
 END
 END vccd_1p0.gds1149
 PIN vccd_1p0.gds1150
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.89 25.8165 39.93 26.0165 ;
 END
 END vccd_1p0.gds1150
 PIN vccd_1p0.gds1151
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 39.218 25.8165 39.258 26.0165 ;
 END
 END vccd_1p0.gds1151
 PIN vccd_1p0.gds1152
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 38.546 25.8165 38.586 26.0165 ;
 END
 END vccd_1p0.gds1152
 PIN vccd_1p0.gds1153
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.874 25.8165 37.914 26.0165 ;
 END
 END vccd_1p0.gds1153
 PIN vccd_1p0.gds1154
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 37.202 25.8165 37.242 26.0165 ;
 END
 END vccd_1p0.gds1154
 PIN vccd_1p0.gds1155
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 36.53 25.8165 36.57 26.0165 ;
 END
 END vccd_1p0.gds1155
 PIN vccd_1p0.gds1156
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.858 25.8165 35.898 26.0165 ;
 END
 END vccd_1p0.gds1156
 PIN vccd_1p0.gds1157
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 40.124 28.1455 40.18 28.3455 ;
 RECT 39.62 28.1755 39.676 28.3755 ;
 RECT 39.452 28.1455 39.508 28.3455 ;
 RECT 39.956 28.044 40.012 28.244 ;
 RECT 38.948 28.1755 39.004 28.3755 ;
 RECT 38.78 28.1455 38.836 28.3455 ;
 RECT 39.284 28.044 39.34 28.244 ;
 RECT 38.276 28.1755 38.332 28.3755 ;
 RECT 38.108 28.1455 38.164 28.3455 ;
 RECT 38.612 28.044 38.668 28.244 ;
 RECT 37.604 28.1755 37.66 28.3755 ;
 RECT 37.436 28.1455 37.492 28.3455 ;
 RECT 37.94 28.044 37.996 28.244 ;
 RECT 36.932 28.1755 36.988 28.3755 ;
 RECT 36.764 28.1455 36.82 28.3455 ;
 RECT 37.268 28.044 37.324 28.244 ;
 RECT 36.26 28.1755 36.316 28.3755 ;
 RECT 36.092 28.1455 36.148 28.3455 ;
 RECT 36.596 28.044 36.652 28.244 ;
 RECT 35.588 28.1755 35.644 28.3755 ;
 RECT 35.252 28.044 35.308 28.244 ;
 RECT 35.42 28.1455 35.476 28.3455 ;
 RECT 35.924 28.044 35.98 28.244 ;
 END
 END vccd_1p0.gds1157
 PIN vccd_1p0.gds1158
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.574 27.6555 44.634 27.8555 ;
 END
 END vccd_1p0.gds1158
 PIN vccd_1p0.gds1159
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.91 27.624 44.97 27.824 ;
 END
 END vccd_1p0.gds1159
 PIN vccd_1p0.gds1160
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.902 27.6555 43.962 27.8555 ;
 END
 END vccd_1p0.gds1160
 PIN vccd_1p0.gds1161
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.238 27.624 44.298 27.824 ;
 END
 END vccd_1p0.gds1161
 PIN vccd_1p0.gds1162
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.23 27.6555 43.29 27.8555 ;
 END
 END vccd_1p0.gds1162
 PIN vccd_1p0.gds1163
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.566 27.624 43.626 27.824 ;
 END
 END vccd_1p0.gds1163
 PIN vccd_1p0.gds1164
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.558 27.6555 42.618 27.8555 ;
 END
 END vccd_1p0.gds1164
 PIN vccd_1p0.gds1165
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.894 27.624 42.954 27.824 ;
 END
 END vccd_1p0.gds1165
 PIN vccd_1p0.gds1166
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.886 27.6555 41.946 27.8555 ;
 END
 END vccd_1p0.gds1166
 PIN vccd_1p0.gds1167
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.222 27.624 42.282 27.824 ;
 END
 END vccd_1p0.gds1167
 PIN vccd_1p0.gds1168
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.214 27.6555 41.274 27.8555 ;
 END
 END vccd_1p0.gds1168
 PIN vccd_1p0.gds1169
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.55 27.624 41.61 27.824 ;
 END
 END vccd_1p0.gds1169
 PIN vccd_1p0.gds1170
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.458 27.624 40.518 27.824 ;
 END
 END vccd_1p0.gds1170
 PIN vccd_1p0.gds1171
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.014 25.8165 45.054 26.0165 ;
 END
 END vccd_1p0.gds1171
 PIN vccd_1p0.gds1172
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 44.342 25.8165 44.382 26.0165 ;
 END
 END vccd_1p0.gds1172
 PIN vccd_1p0.gds1173
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 43.67 25.8165 43.71 26.0165 ;
 END
 END vccd_1p0.gds1173
 PIN vccd_1p0.gds1174
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.998 25.8165 43.038 26.0165 ;
 END
 END vccd_1p0.gds1174
 PIN vccd_1p0.gds1175
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 42.326 25.8165 42.366 26.0165 ;
 END
 END vccd_1p0.gds1175
 PIN vccd_1p0.gds1176
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 41.654 25.8165 41.694 26.0165 ;
 END
 END vccd_1p0.gds1176
 PIN vccd_1p0.gds1177
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.562 25.858 40.602 26.058 ;
 END
 END vccd_1p0.gds1177
 PIN vccd_1p0.gds1178
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 27.9515 40.894 28.1515 ;
 END
 END vccd_1p0.gds1178
 PIN vccd_1p0.gds1179
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 44.744 28.1755 44.8 28.3755 ;
 RECT 44.576 28.1455 44.632 28.3455 ;
 RECT 45.08 28.044 45.136 28.244 ;
 RECT 44.072 28.1755 44.128 28.3755 ;
 RECT 43.904 28.1455 43.96 28.3455 ;
 RECT 44.408 28.044 44.464 28.244 ;
 RECT 43.4 28.1755 43.456 28.3755 ;
 RECT 43.232 28.1455 43.288 28.3455 ;
 RECT 43.736 28.044 43.792 28.244 ;
 RECT 42.728 28.1755 42.784 28.3755 ;
 RECT 42.56 28.1455 42.616 28.3455 ;
 RECT 43.064 28.044 43.12 28.244 ;
 RECT 42.056 28.1755 42.112 28.3755 ;
 RECT 41.888 28.1455 41.944 28.3455 ;
 RECT 42.392 28.044 42.448 28.244 ;
 RECT 41.384 28.1755 41.44 28.3755 ;
 RECT 41.048 28.044 41.104 28.244 ;
 RECT 41.216 28.1455 41.272 28.3455 ;
 RECT 41.72 28.044 41.776 28.244 ;
 RECT 40.628 28.044 40.684 28.244 ;
 RECT 40.292 28.1755 40.348 28.3755 ;
 RECT 40.88 27.6745 40.936 27.8745 ;
 END
 END vccd_1p0.gds1179
 PIN vccd_1p0.gds1180
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.918 27.6555 45.978 27.8555 ;
 END
 END vccd_1p0.gds1180
 PIN vccd_1p0.gds1181
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.254 27.624 46.314 27.824 ;
 END
 END vccd_1p0.gds1181
 PIN vccd_1p0.gds1182
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.246 27.6555 45.306 27.8555 ;
 END
 END vccd_1p0.gds1182
 PIN vccd_1p0.gds1183
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.582 27.624 45.642 27.824 ;
 END
 END vccd_1p0.gds1183
 PIN vccd_1p0.gds1184
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 45.686 25.8165 45.726 26.0165 ;
 END
 END vccd_1p0.gds1184
 PIN vccd_1p0.gds1185
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 29.584 48.082 29.784 ;
 END
 END vccd_1p0.gds1185
 PIN vccd_1p0.gds1186
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 27.777 48.502 27.977 ;
 END
 END vccd_1p0.gds1186
 PIN vccd_1p0.gds1187
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 29.584 48.502 29.784 ;
 END
 END vccd_1p0.gds1187
 PIN vccd_1p0.gds1188
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 29.516 49.394 29.716 ;
 END
 END vccd_1p0.gds1188
 PIN vccd_1p0.gds1189
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 28.6325 47.842 28.8325 ;
 END
 END vccd_1p0.gds1189
 PIN vccd_1p0.gds1190
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 29.075 47.242 29.275 ;
 END
 END vccd_1p0.gds1190
 PIN vccd_1p0.gds1191
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 28.1475 46.758 28.3475 ;
 END
 END vccd_1p0.gds1191
 PIN vccd_1p0.gds1192
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 27.4215 47.002 27.6215 ;
 END
 END vccd_1p0.gds1192
 PIN vccd_1p0.gds1193
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 25.533 48.082 25.733 ;
 END
 END vccd_1p0.gds1193
 PIN vccd_1p0.gds1194
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 28.351 48.082 28.551 ;
 END
 END vccd_1p0.gds1194
 PIN vccd_1p0.gds1195
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 26.687 49.038 26.887 ;
 END
 END vccd_1p0.gds1195
 PIN vccd_1p0.gds1196
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.358 25.8205 46.398 26.0205 ;
 END
 END vccd_1p0.gds1196
 PIN vccd_1p0.gds1197
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 26.8535 48.846 27.0535 ;
 END
 END vccd_1p0.gds1197
 PIN vccd_1p0.gds1198
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 28.0055 49.602 28.2055 ;
 END
 END vccd_1p0.gds1198
 PIN vccd_1p0.gds1199
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 29.7115 49.038 29.9115 ;
 END
 END vccd_1p0.gds1199
 PIN vccd_1p0.gds1200
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 28.28 49.846 28.48 ;
 END
 END vccd_1p0.gds1200
 PIN vccd_1p0.gds1201
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 27.2115 50.33 27.4115 ;
 END
 END vccd_1p0.gds1201
 PIN vccd_1p0.gds1202
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 46.088 28.1755 46.144 28.3755 ;
 RECT 45.92 28.1455 45.976 28.3455 ;
 RECT 46.424 28.044 46.48 28.244 ;
 RECT 45.416 28.1755 45.472 28.3755 ;
 RECT 45.248 28.1455 45.304 28.3455 ;
 RECT 45.752 28.044 45.808 28.244 ;
 RECT 49.364 27.76 49.42 27.96 ;
 RECT 46.844 27.6745 46.9 27.8745 ;
 RECT 47.348 27.486 47.404 27.686 ;
 RECT 46.676 27.76 46.732 27.96 ;
 RECT 49.196 27.76 49.252 27.96 ;
 RECT 49.028 27.854 49.084 28.054 ;
 RECT 48.86 27.6745 48.916 27.8745 ;
 RECT 48.692 27.6745 48.748 27.8745 ;
 RECT 48.524 27.6745 48.58 27.8745 ;
 RECT 48.356 27.6745 48.412 27.8745 ;
 RECT 48.188 27.76 48.244 27.96 ;
 RECT 48.02 27.854 48.076 28.054 ;
 RECT 47.852 27.6745 47.908 27.8745 ;
 RECT 49.7 27.6745 49.756 27.8745 ;
 RECT 49.532 27.76 49.588 27.96 ;
 END
 END vccd_1p0.gds1202
 PIN vccd_1p0.gds1203
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.158 27.6555 55.218 27.8555 ;
 END
 END vccd_1p0.gds1203
 PIN vccd_1p0.gds1204
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.486 27.6555 54.546 27.8555 ;
 END
 END vccd_1p0.gds1204
 PIN vccd_1p0.gds1205
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.822 27.624 54.882 27.824 ;
 END
 END vccd_1p0.gds1205
 PIN vccd_1p0.gds1206
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.814 27.6555 53.874 27.8555 ;
 END
 END vccd_1p0.gds1206
 PIN vccd_1p0.gds1207
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.15 27.624 54.21 27.824 ;
 END
 END vccd_1p0.gds1207
 PIN vccd_1p0.gds1208
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.142 27.6555 53.202 27.8555 ;
 END
 END vccd_1p0.gds1208
 PIN vccd_1p0.gds1209
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.478 27.624 53.538 27.824 ;
 END
 END vccd_1p0.gds1209
 PIN vccd_1p0.gds1210
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.47 27.5315 52.53 27.7315 ;
 END
 END vccd_1p0.gds1210
 PIN vccd_1p0.gds1211
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.806 27.624 52.866 27.824 ;
 END
 END vccd_1p0.gds1211
 PIN vccd_1p0.gds1212
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.926 25.8165 54.966 26.0165 ;
 END
 END vccd_1p0.gds1212
 PIN vccd_1p0.gds1213
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 54.254 25.8165 54.294 26.0165 ;
 END
 END vccd_1p0.gds1213
 PIN vccd_1p0.gds1214
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 53.582 25.8165 53.622 26.0165 ;
 END
 END vccd_1p0.gds1214
 PIN vccd_1p0.gds1215
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 29.648 50.33 29.848 ;
 END
 END vccd_1p0.gds1215
 PIN vccd_1p0.gds1216
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 25.9095 52.194 26.1095 ;
 END
 END vccd_1p0.gds1216
 PIN vccd_1p0.gds1217
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 25.982 52.066 26.182 ;
 END
 END vccd_1p0.gds1217
 PIN vccd_1p0.gds1218
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 27.5675 51.678 27.7675 ;
 END
 END vccd_1p0.gds1218
 PIN vccd_1p0.gds1219
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 29.679 52.194 29.879 ;
 END
 END vccd_1p0.gds1219
 PIN vccd_1p0.gds1220
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 29.5635 52.066 29.7635 ;
 END
 END vccd_1p0.gds1220
 PIN vccd_1p0.gds1221
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 27.223 51.258 27.423 ;
 END
 END vccd_1p0.gds1221
 PIN vccd_1p0.gds1222
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 29.4455 51.838 29.6455 ;
 END
 END vccd_1p0.gds1222
 PIN vccd_1p0.gds1223
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.438 27.875 50.494 28.075 ;
 END
 END vccd_1p0.gds1223
 PIN vccd_1p0.gds1224
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.91 25.8165 52.95 26.0165 ;
 END
 END vccd_1p0.gds1224
 PIN vccd_1p0.gds1225
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 55.16 28.1455 55.216 28.3455 ;
 RECT 54.656 28.1755 54.712 28.3755 ;
 RECT 54.488 28.1455 54.544 28.3455 ;
 RECT 54.992 28.044 55.048 28.244 ;
 RECT 53.984 28.1755 54.04 28.3755 ;
 RECT 53.816 28.1455 53.872 28.3455 ;
 RECT 54.32 28.044 54.376 28.244 ;
 RECT 53.312 28.1755 53.368 28.3755 ;
 RECT 53.144 28.1455 53.2 28.3455 ;
 RECT 53.648 28.044 53.704 28.244 ;
 RECT 52.64 28.1755 52.696 28.3755 ;
 RECT 52.304 28.044 52.36 28.244 ;
 RECT 52.472 28.1455 52.528 28.3455 ;
 RECT 52.976 28.044 53.032 28.244 ;
 RECT 52.052 27.5775 52.108 27.7775 ;
 RECT 51.884 27.76 51.94 27.96 ;
 RECT 51.716 27.6745 51.772 27.8745 ;
 RECT 51.548 27.6745 51.604 27.8745 ;
 RECT 51.38 27.76 51.436 27.96 ;
 RECT 51.212 27.76 51.268 27.96 ;
 END
 END vccd_1p0.gds1225
 PIN vccd_1p0.gds1226
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.61 27.6555 59.67 27.8555 ;
 END
 END vccd_1p0.gds1226
 PIN vccd_1p0.gds1227
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.946 27.624 60.006 27.824 ;
 END
 END vccd_1p0.gds1227
 PIN vccd_1p0.gds1228
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.938 27.6555 58.998 27.8555 ;
 END
 END vccd_1p0.gds1228
 PIN vccd_1p0.gds1229
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.274 27.624 59.334 27.824 ;
 END
 END vccd_1p0.gds1229
 PIN vccd_1p0.gds1230
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.266 27.6555 58.326 27.8555 ;
 END
 END vccd_1p0.gds1230
 PIN vccd_1p0.gds1231
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.602 27.624 58.662 27.824 ;
 END
 END vccd_1p0.gds1231
 PIN vccd_1p0.gds1232
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.174 27.6555 57.234 27.8555 ;
 END
 END vccd_1p0.gds1232
 PIN vccd_1p0.gds1233
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.51 27.624 57.57 27.824 ;
 END
 END vccd_1p0.gds1233
 PIN vccd_1p0.gds1234
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.502 27.6555 56.562 27.8555 ;
 END
 END vccd_1p0.gds1234
 PIN vccd_1p0.gds1235
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.838 27.624 56.898 27.824 ;
 END
 END vccd_1p0.gds1235
 PIN vccd_1p0.gds1236
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.83 27.6555 55.89 27.8555 ;
 END
 END vccd_1p0.gds1236
 PIN vccd_1p0.gds1237
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.166 27.624 56.226 27.824 ;
 END
 END vccd_1p0.gds1237
 PIN vccd_1p0.gds1238
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.494 27.624 55.554 27.824 ;
 END
 END vccd_1p0.gds1238
 PIN vccd_1p0.gds1239
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.05 25.8165 60.09 26.0165 ;
 END
 END vccd_1p0.gds1239
 PIN vccd_1p0.gds1240
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 59.378 25.8165 59.418 26.0165 ;
 END
 END vccd_1p0.gds1240
 PIN vccd_1p0.gds1241
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.942 25.8165 56.982 26.0165 ;
 END
 END vccd_1p0.gds1241
 PIN vccd_1p0.gds1242
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 56.27 25.8165 56.31 26.0165 ;
 END
 END vccd_1p0.gds1242
 PIN vccd_1p0.gds1243
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 55.598 25.8165 55.638 26.0165 ;
 END
 END vccd_1p0.gds1243
 PIN vccd_1p0.gds1244
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 58.706 25.8165 58.746 26.0165 ;
 END
 END vccd_1p0.gds1244
 PIN vccd_1p0.gds1245
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.614 25.858 57.654 26.058 ;
 END
 END vccd_1p0.gds1245
 PIN vccd_1p0.gds1246
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 27.9515 57.946 28.1515 ;
 END
 END vccd_1p0.gds1246
 PIN vccd_1p0.gds1247
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 59.78 28.1755 59.836 28.3755 ;
 RECT 59.612 28.1455 59.668 28.3455 ;
 RECT 60.116 28.044 60.172 28.244 ;
 RECT 59.108 28.1755 59.164 28.3755 ;
 RECT 58.94 28.1455 58.996 28.3455 ;
 RECT 59.444 28.044 59.5 28.244 ;
 RECT 58.436 28.1755 58.492 28.3755 ;
 RECT 58.1 28.044 58.156 28.244 ;
 RECT 58.268 28.1455 58.324 28.3455 ;
 RECT 58.772 28.044 58.828 28.244 ;
 RECT 57.344 28.1755 57.4 28.3755 ;
 RECT 57.176 28.1455 57.232 28.3455 ;
 RECT 57.68 28.044 57.736 28.244 ;
 RECT 56.672 28.1755 56.728 28.3755 ;
 RECT 56.504 28.1455 56.56 28.3455 ;
 RECT 57.008 28.044 57.064 28.244 ;
 RECT 56 28.1755 56.056 28.3755 ;
 RECT 55.832 28.1455 55.888 28.3455 ;
 RECT 56.336 28.044 56.392 28.244 ;
 RECT 55.328 28.1755 55.384 28.3755 ;
 RECT 55.664 28.044 55.72 28.244 ;
 RECT 57.932 27.6745 57.988 27.8745 ;
 END
 END vccd_1p0.gds1247
 PIN vccd_1p0.gds1248
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.97 27.6555 63.03 27.8555 ;
 END
 END vccd_1p0.gds1248
 PIN vccd_1p0.gds1249
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.306 27.624 63.366 27.824 ;
 END
 END vccd_1p0.gds1249
 PIN vccd_1p0.gds1250
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.298 27.6555 62.358 27.8555 ;
 END
 END vccd_1p0.gds1250
 PIN vccd_1p0.gds1251
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.634 27.624 62.694 27.824 ;
 END
 END vccd_1p0.gds1251
 PIN vccd_1p0.gds1252
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.626 27.6555 61.686 27.8555 ;
 END
 END vccd_1p0.gds1252
 PIN vccd_1p0.gds1253
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.962 27.624 62.022 27.824 ;
 END
 END vccd_1p0.gds1253
 PIN vccd_1p0.gds1254
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.954 27.6555 61.014 27.8555 ;
 END
 END vccd_1p0.gds1254
 PIN vccd_1p0.gds1255
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.29 27.624 61.35 27.824 ;
 END
 END vccd_1p0.gds1255
 PIN vccd_1p0.gds1256
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.282 27.6555 60.342 27.8555 ;
 END
 END vccd_1p0.gds1256
 PIN vccd_1p0.gds1257
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.618 27.624 60.678 27.824 ;
 END
 END vccd_1p0.gds1257
 PIN vccd_1p0.gds1258
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.738 25.8165 62.778 26.0165 ;
 END
 END vccd_1p0.gds1258
 PIN vccd_1p0.gds1259
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 62.066 25.8165 62.106 26.0165 ;
 END
 END vccd_1p0.gds1259
 PIN vccd_1p0.gds1260
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 61.394 25.8165 61.434 26.0165 ;
 END
 END vccd_1p0.gds1260
 PIN vccd_1p0.gds1261
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 60.722 25.8165 60.762 26.0165 ;
 END
 END vccd_1p0.gds1261
 PIN vccd_1p0.gds1262
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 29.584 65.134 29.784 ;
 END
 END vccd_1p0.gds1262
 PIN vccd_1p0.gds1263
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 28.6325 64.894 28.8325 ;
 END
 END vccd_1p0.gds1263
 PIN vccd_1p0.gds1264
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 29.075 64.294 29.275 ;
 END
 END vccd_1p0.gds1264
 PIN vccd_1p0.gds1265
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 28.1475 63.81 28.3475 ;
 END
 END vccd_1p0.gds1265
 PIN vccd_1p0.gds1266
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 27.4215 64.054 27.6215 ;
 END
 END vccd_1p0.gds1266
 PIN vccd_1p0.gds1267
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 25.533 65.134 25.733 ;
 END
 END vccd_1p0.gds1267
 PIN vccd_1p0.gds1268
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 28.351 65.134 28.551 ;
 END
 END vccd_1p0.gds1268
 PIN vccd_1p0.gds1269
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.41 25.8205 63.45 26.0205 ;
 END
 END vccd_1p0.gds1269
 PIN vccd_1p0.gds1270
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 63.14 28.1755 63.196 28.3755 ;
 RECT 62.972 28.1455 63.028 28.3455 ;
 RECT 63.476 28.044 63.532 28.244 ;
 RECT 62.468 28.1755 62.524 28.3755 ;
 RECT 62.3 28.1455 62.356 28.3455 ;
 RECT 62.804 28.044 62.86 28.244 ;
 RECT 61.796 28.1755 61.852 28.3755 ;
 RECT 61.628 28.1455 61.684 28.3455 ;
 RECT 62.132 28.044 62.188 28.244 ;
 RECT 61.124 28.1755 61.18 28.3755 ;
 RECT 60.956 28.1455 61.012 28.3455 ;
 RECT 61.46 28.044 61.516 28.244 ;
 RECT 60.452 28.1755 60.508 28.3755 ;
 RECT 60.788 28.044 60.844 28.244 ;
 RECT 60.284 28.1455 60.34 28.3455 ;
 RECT 63.896 27.6745 63.952 27.8745 ;
 RECT 64.4 27.486 64.456 27.686 ;
 RECT 63.728 27.76 63.784 27.96 ;
 RECT 65.072 27.854 65.128 28.054 ;
 RECT 64.904 27.6745 64.96 27.8745 ;
 END
 END vccd_1p0.gds1270
 PIN vccd_1p0.gds1271
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.194 27.6555 70.254 27.8555 ;
 END
 END vccd_1p0.gds1271
 PIN vccd_1p0.gds1272
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.522 27.5315 69.582 27.7315 ;
 END
 END vccd_1p0.gds1272
 PIN vccd_1p0.gds1273
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.858 27.624 69.918 27.824 ;
 END
 END vccd_1p0.gds1273
 PIN vccd_1p0.gds1274
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 25.9095 69.246 26.1095 ;
 END
 END vccd_1p0.gds1274
 PIN vccd_1p0.gds1275
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 25.982 69.118 26.182 ;
 END
 END vccd_1p0.gds1275
 PIN vccd_1p0.gds1276
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 27.777 65.554 27.977 ;
 END
 END vccd_1p0.gds1276
 PIN vccd_1p0.gds1277
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 29.648 67.382 29.848 ;
 END
 END vccd_1p0.gds1277
 PIN vccd_1p0.gds1278
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 29.584 65.554 29.784 ;
 END
 END vccd_1p0.gds1278
 PIN vccd_1p0.gds1279
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 29.516 66.446 29.716 ;
 END
 END vccd_1p0.gds1279
 PIN vccd_1p0.gds1280
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 26.687 66.09 26.887 ;
 END
 END vccd_1p0.gds1280
 PIN vccd_1p0.gds1281
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 26.8535 65.898 27.0535 ;
 END
 END vccd_1p0.gds1281
 PIN vccd_1p0.gds1282
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 27.5675 68.73 27.7675 ;
 END
 END vccd_1p0.gds1282
 PIN vccd_1p0.gds1283
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 29.679 69.246 29.879 ;
 END
 END vccd_1p0.gds1283
 PIN vccd_1p0.gds1284
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 29.5635 69.118 29.7635 ;
 END
 END vccd_1p0.gds1284
 PIN vccd_1p0.gds1285
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 27.223 68.31 27.423 ;
 END
 END vccd_1p0.gds1285
 PIN vccd_1p0.gds1286
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 28.0055 66.654 28.2055 ;
 END
 END vccd_1p0.gds1286
 PIN vccd_1p0.gds1287
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 29.7115 66.09 29.9115 ;
 END
 END vccd_1p0.gds1287
 PIN vccd_1p0.gds1288
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 29.4455 68.89 29.6455 ;
 END
 END vccd_1p0.gds1288
 PIN vccd_1p0.gds1289
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 28.28 66.898 28.48 ;
 END
 END vccd_1p0.gds1289
 PIN vccd_1p0.gds1290
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.49 27.875 67.546 28.075 ;
 END
 END vccd_1p0.gds1290
 PIN vccd_1p0.gds1291
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 27.2115 67.382 27.4115 ;
 END
 END vccd_1p0.gds1291
 PIN vccd_1p0.gds1292
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.962 25.8165 70.002 26.0165 ;
 END
 END vccd_1p0.gds1292
 PIN vccd_1p0.gds1293
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 70.196 28.1455 70.252 28.3455 ;
 RECT 69.692 28.1755 69.748 28.3755 ;
 RECT 69.356 28.044 69.412 28.244 ;
 RECT 69.524 28.1455 69.58 28.3455 ;
 RECT 70.028 28.044 70.084 28.244 ;
 RECT 66.416 27.76 66.472 27.96 ;
 RECT 66.248 27.76 66.304 27.96 ;
 RECT 66.08 27.854 66.136 28.054 ;
 RECT 65.912 27.6745 65.968 27.8745 ;
 RECT 65.744 27.6745 65.8 27.8745 ;
 RECT 65.576 27.6745 65.632 27.8745 ;
 RECT 65.408 27.6745 65.464 27.8745 ;
 RECT 65.24 27.76 65.296 27.96 ;
 RECT 66.752 27.6745 66.808 27.8745 ;
 RECT 66.584 27.76 66.64 27.96 ;
 RECT 69.104 27.5775 69.16 27.7775 ;
 RECT 68.936 27.76 68.992 27.96 ;
 RECT 68.768 27.6745 68.824 27.8745 ;
 RECT 68.6 27.6745 68.656 27.8745 ;
 RECT 68.432 27.76 68.488 27.96 ;
 RECT 68.264 27.76 68.32 27.96 ;
 END
 END vccd_1p0.gds1293
 PIN vccd_1p0.gds1294
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.226 27.6555 74.286 27.8555 ;
 END
 END vccd_1p0.gds1294
 PIN vccd_1p0.gds1295
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.562 27.624 74.622 27.824 ;
 END
 END vccd_1p0.gds1295
 PIN vccd_1p0.gds1296
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.554 27.6555 73.614 27.8555 ;
 END
 END vccd_1p0.gds1296
 PIN vccd_1p0.gds1297
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.89 27.624 73.95 27.824 ;
 END
 END vccd_1p0.gds1297
 PIN vccd_1p0.gds1298
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.882 27.6555 72.942 27.8555 ;
 END
 END vccd_1p0.gds1298
 PIN vccd_1p0.gds1299
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.218 27.624 73.278 27.824 ;
 END
 END vccd_1p0.gds1299
 PIN vccd_1p0.gds1300
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.21 27.6555 72.27 27.8555 ;
 END
 END vccd_1p0.gds1300
 PIN vccd_1p0.gds1301
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.546 27.624 72.606 27.824 ;
 END
 END vccd_1p0.gds1301
 PIN vccd_1p0.gds1302
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.538 27.6555 71.598 27.8555 ;
 END
 END vccd_1p0.gds1302
 PIN vccd_1p0.gds1303
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.874 27.624 71.934 27.824 ;
 END
 END vccd_1p0.gds1303
 PIN vccd_1p0.gds1304
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.866 27.6555 70.926 27.8555 ;
 END
 END vccd_1p0.gds1304
 PIN vccd_1p0.gds1305
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.202 27.624 71.262 27.824 ;
 END
 END vccd_1p0.gds1305
 PIN vccd_1p0.gds1306
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.53 27.624 70.59 27.824 ;
 END
 END vccd_1p0.gds1306
 PIN vccd_1p0.gds1307
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 74.666 25.858 74.706 26.058 ;
 END
 END vccd_1p0.gds1307
 PIN vccd_1p0.gds1308
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.994 25.8165 74.034 26.0165 ;
 END
 END vccd_1p0.gds1308
 PIN vccd_1p0.gds1309
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 73.322 25.8165 73.362 26.0165 ;
 END
 END vccd_1p0.gds1309
 PIN vccd_1p0.gds1310
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 72.65 25.8165 72.69 26.0165 ;
 END
 END vccd_1p0.gds1310
 PIN vccd_1p0.gds1311
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.978 25.8165 72.018 26.0165 ;
 END
 END vccd_1p0.gds1311
 PIN vccd_1p0.gds1312
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 71.306 25.8165 71.346 26.0165 ;
 END
 END vccd_1p0.gds1312
 PIN vccd_1p0.gds1313
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 70.634 25.8165 70.674 26.0165 ;
 END
 END vccd_1p0.gds1313
 PIN vccd_1p0.gds1314
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 74.396 28.1755 74.452 28.3755 ;
 RECT 74.228 28.1455 74.284 28.3455 ;
 RECT 74.732 28.044 74.788 28.244 ;
 RECT 73.724 28.1755 73.78 28.3755 ;
 RECT 73.556 28.1455 73.612 28.3455 ;
 RECT 74.06 28.044 74.116 28.244 ;
 RECT 73.052 28.1755 73.108 28.3755 ;
 RECT 72.884 28.1455 72.94 28.3455 ;
 RECT 73.388 28.044 73.444 28.244 ;
 RECT 72.38 28.1755 72.436 28.3755 ;
 RECT 72.212 28.1455 72.268 28.3455 ;
 RECT 72.716 28.044 72.772 28.244 ;
 RECT 71.708 28.1755 71.764 28.3755 ;
 RECT 71.54 28.1455 71.596 28.3455 ;
 RECT 72.044 28.044 72.1 28.244 ;
 RECT 71.036 28.1755 71.092 28.3755 ;
 RECT 70.868 28.1455 70.924 28.3455 ;
 RECT 71.372 28.044 71.428 28.244 ;
 RECT 70.364 28.1755 70.42 28.3755 ;
 RECT 70.7 28.044 70.756 28.244 ;
 END
 END vccd_1p0.gds1314
 PIN vccd_1p0.gds1315
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 33.218 0.43 33.418 ;
 END
 END vccd_1p0.gds1315
 PIN vccd_1p0.gds1316
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 31.091 4.738 31.291 ;
 END
 END vccd_1p0.gds1316
 PIN vccd_1p0.gds1317
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 35.4195 5.202 35.6195 ;
 END
 END vccd_1p0.gds1317
 PIN vccd_1p0.gds1318
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 34.277 1.542 34.477 ;
 END
 END vccd_1p0.gds1318
 PIN vccd_1p0.gds1319
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 34.1595 5.202 34.3595 ;
 END
 END vccd_1p0.gds1319
 PIN vccd_1p0.gds1320
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 33.017 1.542 33.217 ;
 END
 END vccd_1p0.gds1320
 PIN vccd_1p0.gds1321
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 32.8995 5.202 33.0995 ;
 END
 END vccd_1p0.gds1321
 PIN vccd_1p0.gds1322
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 31.757 1.542 31.957 ;
 END
 END vccd_1p0.gds1322
 PIN vccd_1p0.gds1323
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 31.6395 5.202 31.8395 ;
 END
 END vccd_1p0.gds1323
 PIN vccd_1p0.gds1324
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 30.497 1.542 30.697 ;
 END
 END vccd_1p0.gds1324
 PIN vccd_1p0.gds1325
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 33.362 0.548 33.562 ;
 END
 END vccd_1p0.gds1325
 PIN vccd_1p0.gds1326
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 34.466 1.782 34.666 ;
 END
 END vccd_1p0.gds1326
 PIN vccd_1p0.gds1327
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 33.007 0.858 33.207 ;
 END
 END vccd_1p0.gds1327
 PIN vccd_1p0.gds1328
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 33.212 1.362 33.412 ;
 END
 END vccd_1p0.gds1328
 PIN vccd_1p0.gds1329
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 33.101 1.218 33.301 ;
 END
 END vccd_1p0.gds1329
 PIN vccd_1p0.gds1330
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 33.0635 1.09 33.2635 ;
 END
 END vccd_1p0.gds1330
 PIN vccd_1p0.gds1331
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 35.2245 2.202 35.4245 ;
 END
 END vccd_1p0.gds1331
 PIN vccd_1p0.gds1332
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 32.949 2.622 33.149 ;
 END
 END vccd_1p0.gds1332
 PIN vccd_1p0.gds1333
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 35.4385 2.462 35.6385 ;
 END
 END vccd_1p0.gds1333
 PIN vccd_1p0.gds1334
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 33.0055 3.042 33.2055 ;
 END
 END vccd_1p0.gds1334
 PIN vccd_1p0.gds1335
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 32.641 1.962 32.841 ;
 END
 END vccd_1p0.gds1335
 PIN vccd_1p0.gds1336
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 33.008 2.882 33.208 ;
 END
 END vccd_1p0.gds1336
 PIN vccd_1p0.gds1337
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 33.094 3.39 33.294 ;
 END
 END vccd_1p0.gds1337
 PIN vccd_1p0.gds1338
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 32.92 3.262 33.12 ;
 END
 END vccd_1p0.gds1338
 PIN vccd_1p0.gds1339
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 31.0705 3.666 31.2705 ;
 END
 END vccd_1p0.gds1339
 PIN vccd_1p0.gds1340
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 30.66 4.066 30.86 ;
 END
 END vccd_1p0.gds1340
 PIN vccd_1p0.gds1341
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 31.748 4.258 31.948 ;
 END
 END vccd_1p0.gds1341
 PIN vccd_1p0.gds1342
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 32.9165 3.858 33.1165 ;
 END
 END vccd_1p0.gds1342
 PIN vccd_1p0.gds1343
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 33.102 4.546 33.302 ;
 END
 END vccd_1p0.gds1343
 PIN vccd_1p0.gds1344
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 32.926 5.01 33.126 ;
 END
 END vccd_1p0.gds1344
 PIN vccd_1p0.gds1345
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 4.34 30.712 4.396 30.912 ;
 RECT 4.76 30.688 4.816 30.888 ;
 RECT 5.096 30.712 5.152 30.912 ;
 RECT 4.34 31.972 4.396 32.172 ;
 RECT 4.76 31.948 4.816 32.148 ;
 RECT 5.096 31.972 5.152 32.172 ;
 RECT 4.34 33.232 4.396 33.432 ;
 RECT 4.76 33.208 4.816 33.408 ;
 RECT 5.096 33.232 5.152 33.432 ;
 RECT 4.34 34.492 4.396 34.692 ;
 RECT 4.76 34.468 4.816 34.668 ;
 RECT 5.096 34.492 5.152 34.692 ;
 RECT 3.584 34.3035 3.64 34.5035 ;
 RECT 4.172 34.3895 4.228 34.5895 ;
 RECT 4.928 34.346 4.984 34.546 ;
 RECT 3.584 33.0435 3.64 33.2435 ;
 RECT 4.172 33.1295 4.228 33.3295 ;
 RECT 4.928 33.086 4.984 33.286 ;
 RECT 3.584 31.7835 3.64 31.9835 ;
 RECT 4.172 31.8695 4.228 32.0695 ;
 RECT 4.928 31.826 4.984 32.026 ;
 RECT 3.584 30.5235 3.64 30.7235 ;
 RECT 4.172 30.6095 4.228 30.8095 ;
 RECT 4.928 30.566 4.984 30.766 ;
 END
 END vccd_1p0.gds1345
 PIN vccd_1p0.gds1346
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 32.9165 6.838 33.1165 ;
 END
 END vccd_1p0.gds1346
 PIN vccd_1p0.gds1347
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 33.2335 5.602 33.4335 ;
 END
 END vccd_1p0.gds1347
 PIN vccd_1p0.gds1348
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 31.027 5.41 31.227 ;
 END
 END vccd_1p0.gds1348
 PIN vccd_1p0.gds1349
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 35.024 5.922 35.224 ;
 END
 END vccd_1p0.gds1349
 PIN vccd_1p0.gds1350
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.754 31.2965 5.794 31.4965 ;
 END
 END vccd_1p0.gds1350
 PIN vccd_1p0.gds1351
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 34.133 6.306 34.333 ;
 END
 END vccd_1p0.gds1351
 PIN vccd_1p0.gds1352
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 32.987 6.582 33.187 ;
 END
 END vccd_1p0.gds1352
 PIN vccd_1p0.gds1353
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.6 34.3895 5.656 34.5895 ;
 RECT 5.264 34.3895 5.32 34.5895 ;
 RECT 5.432 34.3035 5.488 34.5035 ;
 RECT 5.936 34.3035 5.992 34.5035 ;
 RECT 5.768 34.3035 5.824 34.5035 ;
 RECT 6.44 34.318 6.496 34.518 ;
 RECT 6.272 34.3035 6.328 34.5035 ;
 RECT 6.104 34.492 6.16 34.692 ;
 RECT 5.6 33.1295 5.656 33.3295 ;
 RECT 5.264 33.1295 5.32 33.3295 ;
 RECT 5.432 33.0435 5.488 33.2435 ;
 RECT 5.936 33.0435 5.992 33.2435 ;
 RECT 5.768 33.0435 5.824 33.2435 ;
 RECT 6.44 33.058 6.496 33.258 ;
 RECT 6.272 33.0435 6.328 33.2435 ;
 RECT 6.104 33.232 6.16 33.432 ;
 RECT 5.6 31.8695 5.656 32.0695 ;
 RECT 5.264 31.8695 5.32 32.0695 ;
 RECT 5.432 31.7835 5.488 31.9835 ;
 RECT 5.936 31.7835 5.992 31.9835 ;
 RECT 5.768 31.7835 5.824 31.9835 ;
 RECT 6.44 31.798 6.496 31.998 ;
 RECT 6.272 31.7835 6.328 31.9835 ;
 RECT 6.104 31.972 6.16 32.172 ;
 RECT 5.6 30.6095 5.656 30.8095 ;
 RECT 5.264 30.6095 5.32 30.8095 ;
 RECT 5.432 30.5235 5.488 30.7235 ;
 RECT 5.936 30.5235 5.992 30.7235 ;
 RECT 5.768 30.5235 5.824 30.7235 ;
 RECT 6.44 30.538 6.496 30.738 ;
 RECT 6.272 30.5235 6.328 30.7235 ;
 RECT 6.104 30.712 6.16 30.912 ;
 END
 END vccd_1p0.gds1353
 PIN vccd_1p0.gds1354
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 30.844 13.978 31.044 ;
 END
 END vccd_1p0.gds1354
 PIN vccd_1p0.gds1355
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 33.364 13.978 33.564 ;
 END
 END vccd_1p0.gds1355
 PIN vccd_1p0.gds1356
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 32.104 13.978 32.304 ;
 END
 END vccd_1p0.gds1356
 PIN vccd_1p0.gds1357
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 34.624 13.978 34.824 ;
 END
 END vccd_1p0.gds1357
 PIN vccd_1p0.gds1358
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 34.624 14.398 34.824 ;
 END
 END vccd_1p0.gds1358
 PIN vccd_1p0.gds1359
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 34.7515 14.934 34.9515 ;
 END
 END vccd_1p0.gds1359
 PIN vccd_1p0.gds1360
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 33.364 14.398 33.564 ;
 END
 END vccd_1p0.gds1360
 PIN vccd_1p0.gds1361
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 33.4915 14.934 33.6915 ;
 END
 END vccd_1p0.gds1361
 PIN vccd_1p0.gds1362
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 32.104 14.398 32.304 ;
 END
 END vccd_1p0.gds1362
 PIN vccd_1p0.gds1363
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 32.2315 14.934 32.4315 ;
 END
 END vccd_1p0.gds1363
 PIN vccd_1p0.gds1364
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 33.984 13.738 34.184 ;
 END
 END vccd_1p0.gds1364
 PIN vccd_1p0.gds1365
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 34.2715 13.138 34.4715 ;
 END
 END vccd_1p0.gds1365
 PIN vccd_1p0.gds1366
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 32.756 12.898 32.956 ;
 END
 END vccd_1p0.gds1366
 PIN vccd_1p0.gds1367
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 33.55 12.654 33.75 ;
 END
 END vccd_1p0.gds1367
 PIN vccd_1p0.gds1368
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 31.0565 12.526 31.2565 ;
 END
 END vccd_1p0.gds1368
 PIN vccd_1p0.gds1369
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 30.844 14.398 31.044 ;
 END
 END vccd_1p0.gds1369
 PIN vccd_1p0.gds1370
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 30.9715 14.934 31.1715 ;
 END
 END vccd_1p0.gds1370
 PIN vccd_1p0.gds1371
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 31.926 14.742 32.126 ;
 END
 END vccd_1p0.gds1371
 PIN vccd_1p0.gds1372
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 30.908 16.226 31.108 ;
 END
 END vccd_1p0.gds1372
 PIN vccd_1p0.gds1373
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 34.688 16.226 34.888 ;
 END
 END vccd_1p0.gds1373
 PIN vccd_1p0.gds1374
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 33.428 16.226 33.628 ;
 END
 END vccd_1p0.gds1374
 PIN vccd_1p0.gds1375
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 32.168 16.226 32.368 ;
 END
 END vccd_1p0.gds1375
 PIN vccd_1p0.gds1376
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 33.798 15.742 33.998 ;
 END
 END vccd_1p0.gds1376
 PIN vccd_1p0.gds1377
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 34.866 15.29 35.066 ;
 END
 END vccd_1p0.gds1377
 PIN vccd_1p0.gds1378
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 32.717 17.574 32.917 ;
 END
 END vccd_1p0.gds1378
 PIN vccd_1p0.gds1379
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 34.6985 18.09 34.8985 ;
 END
 END vccd_1p0.gds1379
 PIN vccd_1p0.gds1380
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 34.81 17.962 35.01 ;
 END
 END vccd_1p0.gds1380
 PIN vccd_1p0.gds1381
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 34.5365 17.734 34.7365 ;
 END
 END vccd_1p0.gds1381
 PIN vccd_1p0.gds1382
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 33.483 15.498 33.683 ;
 END
 END vccd_1p0.gds1382
 PIN vccd_1p0.gds1383
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 32.0135 17.154 32.2135 ;
 END
 END vccd_1p0.gds1383
 PIN vccd_1p0.gds1384
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 32.9875 23.842 33.1875 ;
 END
 END vccd_1p0.gds1384
 PIN vccd_1p0.gds1385
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 33.55 29.706 33.75 ;
 END
 END vccd_1p0.gds1385
 PIN vccd_1p0.gds1386
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 31.0565 29.578 31.2565 ;
 END
 END vccd_1p0.gds1386
 PIN vccd_1p0.gds1387
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 32.756 29.95 32.956 ;
 END
 END vccd_1p0.gds1387
 PIN vccd_1p0.gds1388
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 30.844 31.03 31.044 ;
 END
 END vccd_1p0.gds1388
 PIN vccd_1p0.gds1389
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 34.624 31.03 34.824 ;
 END
 END vccd_1p0.gds1389
 PIN vccd_1p0.gds1390
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 34.688 33.278 34.888 ;
 END
 END vccd_1p0.gds1390
 PIN vccd_1p0.gds1391
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 34.624 31.45 34.824 ;
 END
 END vccd_1p0.gds1391
 PIN vccd_1p0.gds1392
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 34.7515 31.986 34.9515 ;
 END
 END vccd_1p0.gds1392
 PIN vccd_1p0.gds1393
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 33.428 33.278 33.628 ;
 END
 END vccd_1p0.gds1393
 PIN vccd_1p0.gds1394
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 33.364 31.45 33.564 ;
 END
 END vccd_1p0.gds1394
 PIN vccd_1p0.gds1395
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 33.4915 31.986 33.6915 ;
 END
 END vccd_1p0.gds1395
 PIN vccd_1p0.gds1396
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 32.168 33.278 32.368 ;
 END
 END vccd_1p0.gds1396
 PIN vccd_1p0.gds1397
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 32.104 31.45 32.304 ;
 END
 END vccd_1p0.gds1397
 PIN vccd_1p0.gds1398
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 32.2315 31.986 32.4315 ;
 END
 END vccd_1p0.gds1398
 PIN vccd_1p0.gds1399
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 30.908 33.278 31.108 ;
 END
 END vccd_1p0.gds1399
 PIN vccd_1p0.gds1400
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 30.844 31.45 31.044 ;
 END
 END vccd_1p0.gds1400
 PIN vccd_1p0.gds1401
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 30.9715 31.986 31.1715 ;
 END
 END vccd_1p0.gds1401
 PIN vccd_1p0.gds1402
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 34.866 32.342 35.066 ;
 END
 END vccd_1p0.gds1402
 PIN vccd_1p0.gds1403
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 33.364 31.03 33.564 ;
 END
 END vccd_1p0.gds1403
 PIN vccd_1p0.gds1404
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 32.104 31.03 32.304 ;
 END
 END vccd_1p0.gds1404
 PIN vccd_1p0.gds1405
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 33.984 30.79 34.184 ;
 END
 END vccd_1p0.gds1405
 PIN vccd_1p0.gds1406
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 34.2715 30.19 34.4715 ;
 END
 END vccd_1p0.gds1406
 PIN vccd_1p0.gds1407
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 31.926 31.794 32.126 ;
 END
 END vccd_1p0.gds1407
 PIN vccd_1p0.gds1408
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 32.717 34.626 32.917 ;
 END
 END vccd_1p0.gds1408
 PIN vccd_1p0.gds1409
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 34.6985 35.142 34.8985 ;
 END
 END vccd_1p0.gds1409
 PIN vccd_1p0.gds1410
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 34.81 35.014 35.01 ;
 END
 END vccd_1p0.gds1410
 PIN vccd_1p0.gds1411
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 32.0135 34.206 32.2135 ;
 END
 END vccd_1p0.gds1411
 PIN vccd_1p0.gds1412
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 33.483 32.55 33.683 ;
 END
 END vccd_1p0.gds1412
 PIN vccd_1p0.gds1413
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 34.5365 34.786 34.7365 ;
 END
 END vccd_1p0.gds1413
 PIN vccd_1p0.gds1414
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 33.798 32.794 33.998 ;
 END
 END vccd_1p0.gds1414
 PIN vccd_1p0.gds1415
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 32.9875 40.894 33.1875 ;
 END
 END vccd_1p0.gds1415
 PIN vccd_1p0.gds1416
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 30.844 48.082 31.044 ;
 END
 END vccd_1p0.gds1416
 PIN vccd_1p0.gds1417
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 32.104 48.082 32.304 ;
 END
 END vccd_1p0.gds1417
 PIN vccd_1p0.gds1418
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 34.624 48.502 34.824 ;
 END
 END vccd_1p0.gds1418
 PIN vccd_1p0.gds1419
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 34.7515 49.038 34.9515 ;
 END
 END vccd_1p0.gds1419
 PIN vccd_1p0.gds1420
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 33.364 48.502 33.564 ;
 END
 END vccd_1p0.gds1420
 PIN vccd_1p0.gds1421
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 33.4915 49.038 33.6915 ;
 END
 END vccd_1p0.gds1421
 PIN vccd_1p0.gds1422
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 32.104 48.502 32.304 ;
 END
 END vccd_1p0.gds1422
 PIN vccd_1p0.gds1423
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 32.2315 49.038 32.4315 ;
 END
 END vccd_1p0.gds1423
 PIN vccd_1p0.gds1424
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 30.844 48.502 31.044 ;
 END
 END vccd_1p0.gds1424
 PIN vccd_1p0.gds1425
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 30.9715 49.038 31.1715 ;
 END
 END vccd_1p0.gds1425
 PIN vccd_1p0.gds1426
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 34.866 49.394 35.066 ;
 END
 END vccd_1p0.gds1426
 PIN vccd_1p0.gds1427
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 34.624 48.082 34.824 ;
 END
 END vccd_1p0.gds1427
 PIN vccd_1p0.gds1428
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 33.364 48.082 33.564 ;
 END
 END vccd_1p0.gds1428
 PIN vccd_1p0.gds1429
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 33.984 47.842 34.184 ;
 END
 END vccd_1p0.gds1429
 PIN vccd_1p0.gds1430
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 34.2715 47.242 34.4715 ;
 END
 END vccd_1p0.gds1430
 PIN vccd_1p0.gds1431
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 33.55 46.758 33.75 ;
 END
 END vccd_1p0.gds1431
 PIN vccd_1p0.gds1432
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 31.0565 46.63 31.2565 ;
 END
 END vccd_1p0.gds1432
 PIN vccd_1p0.gds1433
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 32.756 47.002 32.956 ;
 END
 END vccd_1p0.gds1433
 PIN vccd_1p0.gds1434
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 31.926 48.846 32.126 ;
 END
 END vccd_1p0.gds1434
 PIN vccd_1p0.gds1435
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 33.483 49.602 33.683 ;
 END
 END vccd_1p0.gds1435
 PIN vccd_1p0.gds1436
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 33.798 49.846 33.998 ;
 END
 END vccd_1p0.gds1436
 PIN vccd_1p0.gds1437
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 34.688 50.33 34.888 ;
 END
 END vccd_1p0.gds1437
 PIN vccd_1p0.gds1438
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 33.428 50.33 33.628 ;
 END
 END vccd_1p0.gds1438
 PIN vccd_1p0.gds1439
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 32.168 50.33 32.368 ;
 END
 END vccd_1p0.gds1439
 PIN vccd_1p0.gds1440
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 30.908 50.33 31.108 ;
 END
 END vccd_1p0.gds1440
 PIN vccd_1p0.gds1441
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 32.717 51.678 32.917 ;
 END
 END vccd_1p0.gds1441
 PIN vccd_1p0.gds1442
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 34.6985 52.194 34.8985 ;
 END
 END vccd_1p0.gds1442
 PIN vccd_1p0.gds1443
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 34.81 52.066 35.01 ;
 END
 END vccd_1p0.gds1443
 PIN vccd_1p0.gds1444
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 32.0135 51.258 32.2135 ;
 END
 END vccd_1p0.gds1444
 PIN vccd_1p0.gds1445
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 34.5365 51.838 34.7365 ;
 END
 END vccd_1p0.gds1445
 PIN vccd_1p0.gds1446
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 32.9875 57.946 33.1875 ;
 END
 END vccd_1p0.gds1446
 PIN vccd_1p0.gds1447
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 30.844 65.134 31.044 ;
 END
 END vccd_1p0.gds1447
 PIN vccd_1p0.gds1448
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 32.104 65.134 32.304 ;
 END
 END vccd_1p0.gds1448
 PIN vccd_1p0.gds1449
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 34.624 65.134 34.824 ;
 END
 END vccd_1p0.gds1449
 PIN vccd_1p0.gds1450
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 33.364 65.134 33.564 ;
 END
 END vccd_1p0.gds1450
 PIN vccd_1p0.gds1451
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 33.984 64.894 34.184 ;
 END
 END vccd_1p0.gds1451
 PIN vccd_1p0.gds1452
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 34.2715 64.294 34.4715 ;
 END
 END vccd_1p0.gds1452
 PIN vccd_1p0.gds1453
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 33.55 63.81 33.75 ;
 END
 END vccd_1p0.gds1453
 PIN vccd_1p0.gds1454
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 31.0565 63.682 31.2565 ;
 END
 END vccd_1p0.gds1454
 PIN vccd_1p0.gds1455
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 32.756 64.054 32.956 ;
 END
 END vccd_1p0.gds1455
 PIN vccd_1p0.gds1456
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 34.688 67.382 34.888 ;
 END
 END vccd_1p0.gds1456
 PIN vccd_1p0.gds1457
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 34.624 65.554 34.824 ;
 END
 END vccd_1p0.gds1457
 PIN vccd_1p0.gds1458
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 34.7515 66.09 34.9515 ;
 END
 END vccd_1p0.gds1458
 PIN vccd_1p0.gds1459
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 33.428 67.382 33.628 ;
 END
 END vccd_1p0.gds1459
 PIN vccd_1p0.gds1460
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 33.364 65.554 33.564 ;
 END
 END vccd_1p0.gds1460
 PIN vccd_1p0.gds1461
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 33.4915 66.09 33.6915 ;
 END
 END vccd_1p0.gds1461
 PIN vccd_1p0.gds1462
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 32.168 67.382 32.368 ;
 END
 END vccd_1p0.gds1462
 PIN vccd_1p0.gds1463
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 32.104 65.554 32.304 ;
 END
 END vccd_1p0.gds1463
 PIN vccd_1p0.gds1464
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 32.2315 66.09 32.4315 ;
 END
 END vccd_1p0.gds1464
 PIN vccd_1p0.gds1465
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 30.908 67.382 31.108 ;
 END
 END vccd_1p0.gds1465
 PIN vccd_1p0.gds1466
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 30.844 65.554 31.044 ;
 END
 END vccd_1p0.gds1466
 PIN vccd_1p0.gds1467
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 30.9715 66.09 31.1715 ;
 END
 END vccd_1p0.gds1467
 PIN vccd_1p0.gds1468
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 34.866 66.446 35.066 ;
 END
 END vccd_1p0.gds1468
 PIN vccd_1p0.gds1469
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 31.926 65.898 32.126 ;
 END
 END vccd_1p0.gds1469
 PIN vccd_1p0.gds1470
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 32.717 68.73 32.917 ;
 END
 END vccd_1p0.gds1470
 PIN vccd_1p0.gds1471
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 34.6985 69.246 34.8985 ;
 END
 END vccd_1p0.gds1471
 PIN vccd_1p0.gds1472
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 34.81 69.118 35.01 ;
 END
 END vccd_1p0.gds1472
 PIN vccd_1p0.gds1473
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 32.0135 68.31 32.2135 ;
 END
 END vccd_1p0.gds1473
 PIN vccd_1p0.gds1474
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 33.483 66.654 33.683 ;
 END
 END vccd_1p0.gds1474
 PIN vccd_1p0.gds1475
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 34.5365 68.89 34.7365 ;
 END
 END vccd_1p0.gds1475
 PIN vccd_1p0.gds1476
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 33.798 66.898 33.998 ;
 END
 END vccd_1p0.gds1476
 PIN vccd_1p0.gds1477
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 38.131 0.43 38.331 ;
 END
 END vccd_1p0.gds1477
 PIN vccd_1p0.gds1478
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 36.0715 4.738 36.2715 ;
 END
 END vccd_1p0.gds1478
 PIN vccd_1p0.gds1479
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 39.317 1.542 39.517 ;
 END
 END vccd_1p0.gds1479
 PIN vccd_1p0.gds1480
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 36.797 1.542 36.997 ;
 END
 END vccd_1p0.gds1480
 PIN vccd_1p0.gds1481
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 35.537 1.542 35.737 ;
 END
 END vccd_1p0.gds1481
 PIN vccd_1p0.gds1482
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 38.057 1.542 38.257 ;
 END
 END vccd_1p0.gds1482
 PIN vccd_1p0.gds1483
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 38.243 0.548 38.443 ;
 END
 END vccd_1p0.gds1483
 PIN vccd_1p0.gds1484
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 39.506 1.782 39.706 ;
 END
 END vccd_1p0.gds1484
 PIN vccd_1p0.gds1485
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 38.047 0.858 38.247 ;
 END
 END vccd_1p0.gds1485
 PIN vccd_1p0.gds1486
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 38.252 1.362 38.452 ;
 END
 END vccd_1p0.gds1486
 PIN vccd_1p0.gds1487
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 38.141 1.218 38.341 ;
 END
 END vccd_1p0.gds1487
 PIN vccd_1p0.gds1488
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 38.1035 1.09 38.3035 ;
 END
 END vccd_1p0.gds1488
 PIN vccd_1p0.gds1489
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 40.2645 2.202 40.4645 ;
 END
 END vccd_1p0.gds1489
 PIN vccd_1p0.gds1490
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 37.989 2.622 38.189 ;
 END
 END vccd_1p0.gds1490
 PIN vccd_1p0.gds1491
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 40.4085 2.462 40.6085 ;
 END
 END vccd_1p0.gds1491
 PIN vccd_1p0.gds1492
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 38.0455 3.042 38.2455 ;
 END
 END vccd_1p0.gds1492
 PIN vccd_1p0.gds1493
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 37.9395 5.202 38.1395 ;
 END
 END vccd_1p0.gds1493
 PIN vccd_1p0.gds1494
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 39.1995 5.202 39.3995 ;
 END
 END vccd_1p0.gds1494
 PIN vccd_1p0.gds1495
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 37.681 1.962 37.881 ;
 END
 END vccd_1p0.gds1495
 PIN vccd_1p0.gds1496
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 38.048 2.882 38.248 ;
 END
 END vccd_1p0.gds1496
 PIN vccd_1p0.gds1497
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 38.134 3.39 38.334 ;
 END
 END vccd_1p0.gds1497
 PIN vccd_1p0.gds1498
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 37.96 3.262 38.16 ;
 END
 END vccd_1p0.gds1498
 PIN vccd_1p0.gds1499
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 36.6795 5.202 36.8795 ;
 END
 END vccd_1p0.gds1499
 PIN vccd_1p0.gds1500
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 36.0065 3.666 36.2065 ;
 END
 END vccd_1p0.gds1500
 PIN vccd_1p0.gds1501
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 35.6165 4.066 35.8165 ;
 END
 END vccd_1p0.gds1501
 PIN vccd_1p0.gds1502
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 36.788 4.258 36.988 ;
 END
 END vccd_1p0.gds1502
 PIN vccd_1p0.gds1503
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 37.9565 3.858 38.1565 ;
 END
 END vccd_1p0.gds1503
 PIN vccd_1p0.gds1504
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 38.07 4.546 38.27 ;
 END
 END vccd_1p0.gds1504
 PIN vccd_1p0.gds1505
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 37.966 5.01 38.166 ;
 END
 END vccd_1p0.gds1505
 PIN vccd_1p0.gds1506
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 4.34 35.752 4.396 35.952 ;
 RECT 4.76 35.728 4.816 35.928 ;
 RECT 5.096 35.752 5.152 35.952 ;
 RECT 4.34 37.012 4.396 37.212 ;
 RECT 4.76 36.988 4.816 37.188 ;
 RECT 5.096 37.012 5.152 37.212 ;
 RECT 4.34 38.272 4.396 38.472 ;
 RECT 4.76 38.248 4.816 38.448 ;
 RECT 5.096 38.272 5.152 38.472 ;
 RECT 4.34 39.532 4.396 39.732 ;
 RECT 4.76 39.508 4.816 39.708 ;
 RECT 5.096 39.532 5.152 39.732 ;
 RECT 3.584 39.3435 3.64 39.5435 ;
 RECT 4.172 39.4295 4.228 39.6295 ;
 RECT 4.928 39.386 4.984 39.586 ;
 RECT 3.584 38.0835 3.64 38.2835 ;
 RECT 4.172 38.1695 4.228 38.3695 ;
 RECT 4.928 38.126 4.984 38.326 ;
 RECT 3.584 36.8235 3.64 37.0235 ;
 RECT 4.172 36.9095 4.228 37.1095 ;
 RECT 4.928 36.866 4.984 37.066 ;
 RECT 3.584 35.5635 3.64 35.7635 ;
 RECT 4.172 35.6495 4.228 35.8495 ;
 RECT 4.928 35.606 4.984 35.806 ;
 END
 END vccd_1p0.gds1506
 PIN vccd_1p0.gds1507
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 37.9565 6.838 38.1565 ;
 END
 END vccd_1p0.gds1507
 PIN vccd_1p0.gds1508
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 38.1135 5.602 38.3135 ;
 END
 END vccd_1p0.gds1508
 PIN vccd_1p0.gds1509
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 35.446 6.05 35.646 ;
 END
 END vccd_1p0.gds1509
 PIN vccd_1p0.gds1510
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 35.9765 5.41 36.1765 ;
 END
 END vccd_1p0.gds1510
 PIN vccd_1p0.gds1511
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 40.064 5.922 40.264 ;
 END
 END vccd_1p0.gds1511
 PIN vccd_1p0.gds1512
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.754 36.3365 5.794 36.5365 ;
 END
 END vccd_1p0.gds1512
 PIN vccd_1p0.gds1513
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 39.173 6.306 39.373 ;
 END
 END vccd_1p0.gds1513
 PIN vccd_1p0.gds1514
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 38.027 6.582 38.227 ;
 END
 END vccd_1p0.gds1514
 PIN vccd_1p0.gds1515
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.6 39.4295 5.656 39.6295 ;
 RECT 5.264 39.4295 5.32 39.6295 ;
 RECT 5.432 39.3435 5.488 39.5435 ;
 RECT 5.936 39.3435 5.992 39.5435 ;
 RECT 5.768 39.3435 5.824 39.5435 ;
 RECT 6.44 39.358 6.496 39.558 ;
 RECT 6.272 39.3435 6.328 39.5435 ;
 RECT 6.104 39.532 6.16 39.732 ;
 RECT 5.6 38.1695 5.656 38.3695 ;
 RECT 5.264 38.1695 5.32 38.3695 ;
 RECT 5.432 38.0835 5.488 38.2835 ;
 RECT 5.936 38.0835 5.992 38.2835 ;
 RECT 5.768 38.0835 5.824 38.2835 ;
 RECT 6.44 38.098 6.496 38.298 ;
 RECT 6.272 38.0835 6.328 38.2835 ;
 RECT 6.104 38.272 6.16 38.472 ;
 RECT 5.6 36.9095 5.656 37.1095 ;
 RECT 5.264 36.9095 5.32 37.1095 ;
 RECT 5.432 36.8235 5.488 37.0235 ;
 RECT 5.936 36.8235 5.992 37.0235 ;
 RECT 5.768 36.8235 5.824 37.0235 ;
 RECT 6.44 36.838 6.496 37.038 ;
 RECT 6.272 36.8235 6.328 37.0235 ;
 RECT 6.104 37.012 6.16 37.212 ;
 RECT 5.6 35.6495 5.656 35.8495 ;
 RECT 5.264 35.6495 5.32 35.8495 ;
 RECT 5.432 35.5635 5.488 35.7635 ;
 RECT 5.936 35.5635 5.992 35.7635 ;
 RECT 5.768 35.5635 5.824 35.7635 ;
 RECT 6.44 35.578 6.496 35.778 ;
 RECT 6.272 35.5635 6.328 35.7635 ;
 RECT 6.104 35.752 6.16 35.952 ;
 END
 END vccd_1p0.gds1515
 PIN vccd_1p0.gds1516
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 35.884 13.978 36.084 ;
 END
 END vccd_1p0.gds1516
 PIN vccd_1p0.gds1517
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 37.144 13.978 37.344 ;
 END
 END vccd_1p0.gds1517
 PIN vccd_1p0.gds1518
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 38.404 13.978 38.604 ;
 END
 END vccd_1p0.gds1518
 PIN vccd_1p0.gds1519
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 39.664 13.978 39.864 ;
 END
 END vccd_1p0.gds1519
 PIN vccd_1p0.gds1520
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 35.884 14.398 36.084 ;
 END
 END vccd_1p0.gds1520
 PIN vccd_1p0.gds1521
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 36.0115 14.934 36.2115 ;
 END
 END vccd_1p0.gds1521
 PIN vccd_1p0.gds1522
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 37.144 14.398 37.344 ;
 END
 END vccd_1p0.gds1522
 PIN vccd_1p0.gds1523
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 37.2715 14.934 37.4715 ;
 END
 END vccd_1p0.gds1523
 PIN vccd_1p0.gds1524
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 38.404 14.398 38.604 ;
 END
 END vccd_1p0.gds1524
 PIN vccd_1p0.gds1525
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 38.5315 14.934 38.7315 ;
 END
 END vccd_1p0.gds1525
 PIN vccd_1p0.gds1526
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 39.664 14.398 39.864 ;
 END
 END vccd_1p0.gds1526
 PIN vccd_1p0.gds1527
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 39.7915 14.934 39.9915 ;
 END
 END vccd_1p0.gds1527
 PIN vccd_1p0.gds1528
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 39.024 13.738 39.224 ;
 END
 END vccd_1p0.gds1528
 PIN vccd_1p0.gds1529
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 39.3115 13.138 39.5115 ;
 END
 END vccd_1p0.gds1529
 PIN vccd_1p0.gds1530
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 37.6725 12.898 37.8725 ;
 END
 END vccd_1p0.gds1530
 PIN vccd_1p0.gds1531
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 38.59 12.654 38.79 ;
 END
 END vccd_1p0.gds1531
 PIN vccd_1p0.gds1532
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 36.028 12.526 36.228 ;
 END
 END vccd_1p0.gds1532
 PIN vccd_1p0.gds1533
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 36.7435 14.742 36.9435 ;
 END
 END vccd_1p0.gds1533
 PIN vccd_1p0.gds1534
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 35.948 16.226 36.148 ;
 END
 END vccd_1p0.gds1534
 PIN vccd_1p0.gds1535
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 37.208 16.226 37.408 ;
 END
 END vccd_1p0.gds1535
 PIN vccd_1p0.gds1536
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 38.468 16.226 38.668 ;
 END
 END vccd_1p0.gds1536
 PIN vccd_1p0.gds1537
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 39.728 16.226 39.928 ;
 END
 END vccd_1p0.gds1537
 PIN vccd_1p0.gds1538
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 38.838 15.742 39.038 ;
 END
 END vccd_1p0.gds1538
 PIN vccd_1p0.gds1539
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 39.906 15.29 40.106 ;
 END
 END vccd_1p0.gds1539
 PIN vccd_1p0.gds1540
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 37.757 17.574 37.957 ;
 END
 END vccd_1p0.gds1540
 PIN vccd_1p0.gds1541
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 39.7385 18.09 39.9385 ;
 END
 END vccd_1p0.gds1541
 PIN vccd_1p0.gds1542
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 39.85 17.962 40.05 ;
 END
 END vccd_1p0.gds1542
 PIN vccd_1p0.gds1543
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 39.5765 17.734 39.7765 ;
 END
 END vccd_1p0.gds1543
 PIN vccd_1p0.gds1544
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 38.523 15.498 38.723 ;
 END
 END vccd_1p0.gds1544
 PIN vccd_1p0.gds1545
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 36.8965 17.154 37.0965 ;
 END
 END vccd_1p0.gds1545
 PIN vccd_1p0.gds1546
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 38.0275 23.842 38.2275 ;
 END
 END vccd_1p0.gds1546
 PIN vccd_1p0.gds1547
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 38.59 29.706 38.79 ;
 END
 END vccd_1p0.gds1547
 PIN vccd_1p0.gds1548
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 36.028 29.578 36.228 ;
 END
 END vccd_1p0.gds1548
 PIN vccd_1p0.gds1549
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 37.6725 29.95 37.8725 ;
 END
 END vccd_1p0.gds1549
 PIN vccd_1p0.gds1550
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 35.884 31.03 36.084 ;
 END
 END vccd_1p0.gds1550
 PIN vccd_1p0.gds1551
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 39.728 33.278 39.928 ;
 END
 END vccd_1p0.gds1551
 PIN vccd_1p0.gds1552
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 39.664 31.45 39.864 ;
 END
 END vccd_1p0.gds1552
 PIN vccd_1p0.gds1553
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 39.7915 31.986 39.9915 ;
 END
 END vccd_1p0.gds1553
 PIN vccd_1p0.gds1554
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 37.208 33.278 37.408 ;
 END
 END vccd_1p0.gds1554
 PIN vccd_1p0.gds1555
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 37.144 31.45 37.344 ;
 END
 END vccd_1p0.gds1555
 PIN vccd_1p0.gds1556
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 37.2715 31.986 37.4715 ;
 END
 END vccd_1p0.gds1556
 PIN vccd_1p0.gds1557
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 35.948 33.278 36.148 ;
 END
 END vccd_1p0.gds1557
 PIN vccd_1p0.gds1558
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 35.884 31.45 36.084 ;
 END
 END vccd_1p0.gds1558
 PIN vccd_1p0.gds1559
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 36.0115 31.986 36.2115 ;
 END
 END vccd_1p0.gds1559
 PIN vccd_1p0.gds1560
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 38.468 33.278 38.668 ;
 END
 END vccd_1p0.gds1560
 PIN vccd_1p0.gds1561
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 38.404 31.45 38.604 ;
 END
 END vccd_1p0.gds1561
 PIN vccd_1p0.gds1562
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 38.5315 31.986 38.7315 ;
 END
 END vccd_1p0.gds1562
 PIN vccd_1p0.gds1563
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 39.906 32.342 40.106 ;
 END
 END vccd_1p0.gds1563
 PIN vccd_1p0.gds1564
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 37.144 31.03 37.344 ;
 END
 END vccd_1p0.gds1564
 PIN vccd_1p0.gds1565
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 38.404 31.03 38.604 ;
 END
 END vccd_1p0.gds1565
 PIN vccd_1p0.gds1566
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 39.664 31.03 39.864 ;
 END
 END vccd_1p0.gds1566
 PIN vccd_1p0.gds1567
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 39.024 30.79 39.224 ;
 END
 END vccd_1p0.gds1567
 PIN vccd_1p0.gds1568
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 39.3115 30.19 39.5115 ;
 END
 END vccd_1p0.gds1568
 PIN vccd_1p0.gds1569
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 36.7435 31.794 36.9435 ;
 END
 END vccd_1p0.gds1569
 PIN vccd_1p0.gds1570
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 37.757 34.626 37.957 ;
 END
 END vccd_1p0.gds1570
 PIN vccd_1p0.gds1571
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 39.7385 35.142 39.9385 ;
 END
 END vccd_1p0.gds1571
 PIN vccd_1p0.gds1572
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 39.85 35.014 40.05 ;
 END
 END vccd_1p0.gds1572
 PIN vccd_1p0.gds1573
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 36.8965 34.206 37.0965 ;
 END
 END vccd_1p0.gds1573
 PIN vccd_1p0.gds1574
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 38.523 32.55 38.723 ;
 END
 END vccd_1p0.gds1574
 PIN vccd_1p0.gds1575
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 39.5765 34.786 39.7765 ;
 END
 END vccd_1p0.gds1575
 PIN vccd_1p0.gds1576
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 38.838 32.794 39.038 ;
 END
 END vccd_1p0.gds1576
 PIN vccd_1p0.gds1577
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 38.0275 40.894 38.2275 ;
 END
 END vccd_1p0.gds1577
 PIN vccd_1p0.gds1578
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 38.404 48.082 38.604 ;
 END
 END vccd_1p0.gds1578
 PIN vccd_1p0.gds1579
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 39.664 48.082 39.864 ;
 END
 END vccd_1p0.gds1579
 PIN vccd_1p0.gds1580
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 37.144 48.082 37.344 ;
 END
 END vccd_1p0.gds1580
 PIN vccd_1p0.gds1581
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 35.884 48.082 36.084 ;
 END
 END vccd_1p0.gds1581
 PIN vccd_1p0.gds1582
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 37.144 48.502 37.344 ;
 END
 END vccd_1p0.gds1582
 PIN vccd_1p0.gds1583
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 37.2715 49.038 37.4715 ;
 END
 END vccd_1p0.gds1583
 PIN vccd_1p0.gds1584
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 38.404 48.502 38.604 ;
 END
 END vccd_1p0.gds1584
 PIN vccd_1p0.gds1585
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 38.5315 49.038 38.7315 ;
 END
 END vccd_1p0.gds1585
 PIN vccd_1p0.gds1586
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 39.664 48.502 39.864 ;
 END
 END vccd_1p0.gds1586
 PIN vccd_1p0.gds1587
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 39.7915 49.038 39.9915 ;
 END
 END vccd_1p0.gds1587
 PIN vccd_1p0.gds1588
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 35.884 48.502 36.084 ;
 END
 END vccd_1p0.gds1588
 PIN vccd_1p0.gds1589
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 36.0115 49.038 36.2115 ;
 END
 END vccd_1p0.gds1589
 PIN vccd_1p0.gds1590
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 39.906 49.394 40.106 ;
 END
 END vccd_1p0.gds1590
 PIN vccd_1p0.gds1591
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 39.024 47.842 39.224 ;
 END
 END vccd_1p0.gds1591
 PIN vccd_1p0.gds1592
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 39.3115 47.242 39.5115 ;
 END
 END vccd_1p0.gds1592
 PIN vccd_1p0.gds1593
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 38.59 46.758 38.79 ;
 END
 END vccd_1p0.gds1593
 PIN vccd_1p0.gds1594
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 36.028 46.63 36.228 ;
 END
 END vccd_1p0.gds1594
 PIN vccd_1p0.gds1595
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 37.6725 47.002 37.8725 ;
 END
 END vccd_1p0.gds1595
 PIN vccd_1p0.gds1596
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 36.7435 48.846 36.9435 ;
 END
 END vccd_1p0.gds1596
 PIN vccd_1p0.gds1597
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 38.523 49.602 38.723 ;
 END
 END vccd_1p0.gds1597
 PIN vccd_1p0.gds1598
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 38.838 49.846 39.038 ;
 END
 END vccd_1p0.gds1598
 PIN vccd_1p0.gds1599
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 37.208 50.33 37.408 ;
 END
 END vccd_1p0.gds1599
 PIN vccd_1p0.gds1600
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 38.468 50.33 38.668 ;
 END
 END vccd_1p0.gds1600
 PIN vccd_1p0.gds1601
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 39.728 50.33 39.928 ;
 END
 END vccd_1p0.gds1601
 PIN vccd_1p0.gds1602
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 35.948 50.33 36.148 ;
 END
 END vccd_1p0.gds1602
 PIN vccd_1p0.gds1603
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 37.757 51.678 37.957 ;
 END
 END vccd_1p0.gds1603
 PIN vccd_1p0.gds1604
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 39.7385 52.194 39.9385 ;
 END
 END vccd_1p0.gds1604
 PIN vccd_1p0.gds1605
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 39.85 52.066 40.05 ;
 END
 END vccd_1p0.gds1605
 PIN vccd_1p0.gds1606
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 36.8965 51.258 37.0965 ;
 END
 END vccd_1p0.gds1606
 PIN vccd_1p0.gds1607
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 39.5765 51.838 39.7765 ;
 END
 END vccd_1p0.gds1607
 PIN vccd_1p0.gds1608
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 38.0275 57.946 38.2275 ;
 END
 END vccd_1p0.gds1608
 PIN vccd_1p0.gds1609
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 35.884 65.134 36.084 ;
 END
 END vccd_1p0.gds1609
 PIN vccd_1p0.gds1610
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 37.144 65.134 37.344 ;
 END
 END vccd_1p0.gds1610
 PIN vccd_1p0.gds1611
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 38.404 65.134 38.604 ;
 END
 END vccd_1p0.gds1611
 PIN vccd_1p0.gds1612
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 39.664 65.134 39.864 ;
 END
 END vccd_1p0.gds1612
 PIN vccd_1p0.gds1613
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 39.024 64.894 39.224 ;
 END
 END vccd_1p0.gds1613
 PIN vccd_1p0.gds1614
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 39.3115 64.294 39.5115 ;
 END
 END vccd_1p0.gds1614
 PIN vccd_1p0.gds1615
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 38.59 63.81 38.79 ;
 END
 END vccd_1p0.gds1615
 PIN vccd_1p0.gds1616
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 36.028 63.682 36.228 ;
 END
 END vccd_1p0.gds1616
 PIN vccd_1p0.gds1617
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 37.6725 64.054 37.8725 ;
 END
 END vccd_1p0.gds1617
 PIN vccd_1p0.gds1618
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 37.208 67.382 37.408 ;
 END
 END vccd_1p0.gds1618
 PIN vccd_1p0.gds1619
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 37.144 65.554 37.344 ;
 END
 END vccd_1p0.gds1619
 PIN vccd_1p0.gds1620
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 37.2715 66.09 37.4715 ;
 END
 END vccd_1p0.gds1620
 PIN vccd_1p0.gds1621
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 38.468 67.382 38.668 ;
 END
 END vccd_1p0.gds1621
 PIN vccd_1p0.gds1622
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 38.404 65.554 38.604 ;
 END
 END vccd_1p0.gds1622
 PIN vccd_1p0.gds1623
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 38.5315 66.09 38.7315 ;
 END
 END vccd_1p0.gds1623
 PIN vccd_1p0.gds1624
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 39.728 67.382 39.928 ;
 END
 END vccd_1p0.gds1624
 PIN vccd_1p0.gds1625
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 39.664 65.554 39.864 ;
 END
 END vccd_1p0.gds1625
 PIN vccd_1p0.gds1626
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 39.7915 66.09 39.9915 ;
 END
 END vccd_1p0.gds1626
 PIN vccd_1p0.gds1627
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 35.948 67.382 36.148 ;
 END
 END vccd_1p0.gds1627
 PIN vccd_1p0.gds1628
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 35.884 65.554 36.084 ;
 END
 END vccd_1p0.gds1628
 PIN vccd_1p0.gds1629
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 36.0115 66.09 36.2115 ;
 END
 END vccd_1p0.gds1629
 PIN vccd_1p0.gds1630
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 39.906 66.446 40.106 ;
 END
 END vccd_1p0.gds1630
 PIN vccd_1p0.gds1631
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 36.7435 65.898 36.9435 ;
 END
 END vccd_1p0.gds1631
 PIN vccd_1p0.gds1632
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 37.757 68.73 37.957 ;
 END
 END vccd_1p0.gds1632
 PIN vccd_1p0.gds1633
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 39.7385 69.246 39.9385 ;
 END
 END vccd_1p0.gds1633
 PIN vccd_1p0.gds1634
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 39.85 69.118 40.05 ;
 END
 END vccd_1p0.gds1634
 PIN vccd_1p0.gds1635
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 36.8965 68.31 37.0965 ;
 END
 END vccd_1p0.gds1635
 PIN vccd_1p0.gds1636
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 38.523 66.654 38.723 ;
 END
 END vccd_1p0.gds1636
 PIN vccd_1p0.gds1637
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 39.5765 68.89 39.7765 ;
 END
 END vccd_1p0.gds1637
 PIN vccd_1p0.gds1638
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 38.838 66.898 39.038 ;
 END
 END vccd_1p0.gds1638
 PIN vccd_1p0.gds1639
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 43.046 0.43 43.246 ;
 END
 END vccd_1p0.gds1639
 PIN vccd_1p0.gds1640
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 40.9845 4.738 41.1845 ;
 END
 END vccd_1p0.gds1640
 PIN vccd_1p0.gds1641
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 40.577 1.542 40.777 ;
 END
 END vccd_1p0.gds1641
 PIN vccd_1p0.gds1642
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 41.837 1.542 42.037 ;
 END
 END vccd_1p0.gds1642
 PIN vccd_1p0.gds1643
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 43.097 1.542 43.297 ;
 END
 END vccd_1p0.gds1643
 PIN vccd_1p0.gds1644
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 42.9795 5.202 43.1795 ;
 END
 END vccd_1p0.gds1644
 PIN vccd_1p0.gds1645
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 44.357 1.542 44.557 ;
 END
 END vccd_1p0.gds1645
 PIN vccd_1p0.gds1646
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 43.283 0.548 43.483 ;
 END
 END vccd_1p0.gds1646
 PIN vccd_1p0.gds1647
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 44.546 1.782 44.746 ;
 END
 END vccd_1p0.gds1647
 PIN vccd_1p0.gds1648
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 43.0055 0.858 43.2055 ;
 END
 END vccd_1p0.gds1648
 PIN vccd_1p0.gds1649
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 43.292 1.362 43.492 ;
 END
 END vccd_1p0.gds1649
 PIN vccd_1p0.gds1650
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 43.181 1.218 43.381 ;
 END
 END vccd_1p0.gds1650
 PIN vccd_1p0.gds1651
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 43.0865 1.09 43.2865 ;
 END
 END vccd_1p0.gds1651
 PIN vccd_1p0.gds1652
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 45.3045 2.202 45.5045 ;
 END
 END vccd_1p0.gds1652
 PIN vccd_1p0.gds1653
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 42.973 2.622 43.173 ;
 END
 END vccd_1p0.gds1653
 PIN vccd_1p0.gds1654
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 45.3785 2.462 45.5785 ;
 END
 END vccd_1p0.gds1654
 PIN vccd_1p0.gds1655
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 44.2395 5.202 44.4395 ;
 END
 END vccd_1p0.gds1655
 PIN vccd_1p0.gds1656
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 41.7195 5.202 41.9195 ;
 END
 END vccd_1p0.gds1656
 PIN vccd_1p0.gds1657
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 43.0855 3.042 43.2855 ;
 END
 END vccd_1p0.gds1657
 PIN vccd_1p0.gds1658
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 40.4595 5.202 40.6595 ;
 END
 END vccd_1p0.gds1658
 PIN vccd_1p0.gds1659
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 42.721 1.962 42.921 ;
 END
 END vccd_1p0.gds1659
 PIN vccd_1p0.gds1660
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 43.088 2.882 43.288 ;
 END
 END vccd_1p0.gds1660
 PIN vccd_1p0.gds1661
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 43.174 3.39 43.374 ;
 END
 END vccd_1p0.gds1661
 PIN vccd_1p0.gds1662
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 43 3.262 43.2 ;
 END
 END vccd_1p0.gds1662
 PIN vccd_1p0.gds1663
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 40.943 3.666 41.143 ;
 END
 END vccd_1p0.gds1663
 PIN vccd_1p0.gds1664
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 40.6565 4.066 40.8565 ;
 END
 END vccd_1p0.gds1664
 PIN vccd_1p0.gds1665
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 41.828 4.258 42.028 ;
 END
 END vccd_1p0.gds1665
 PIN vccd_1p0.gds1666
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 42.9965 3.858 43.1965 ;
 END
 END vccd_1p0.gds1666
 PIN vccd_1p0.gds1667
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 43.042 4.546 43.242 ;
 END
 END vccd_1p0.gds1667
 PIN vccd_1p0.gds1668
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 43.006 5.01 43.206 ;
 END
 END vccd_1p0.gds1668
 PIN vccd_1p0.gds1669
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 4.34 42.052 4.396 42.252 ;
 RECT 4.76 42.028 4.816 42.228 ;
 RECT 5.096 42.052 5.152 42.252 ;
 RECT 4.34 43.312 4.396 43.512 ;
 RECT 4.76 43.288 4.816 43.488 ;
 RECT 5.096 43.312 5.152 43.512 ;
 RECT 4.34 44.572 4.396 44.772 ;
 RECT 4.76 44.548 4.816 44.748 ;
 RECT 5.096 44.572 5.152 44.772 ;
 RECT 3.584 44.3835 3.64 44.5835 ;
 RECT 4.172 44.4695 4.228 44.6695 ;
 RECT 4.928 44.426 4.984 44.626 ;
 RECT 3.584 43.1235 3.64 43.3235 ;
 RECT 4.172 43.2095 4.228 43.4095 ;
 RECT 4.928 43.166 4.984 43.366 ;
 RECT 3.584 41.8635 3.64 42.0635 ;
 RECT 4.172 41.9495 4.228 42.1495 ;
 RECT 4.928 41.906 4.984 42.106 ;
 RECT 4.34 40.792 4.396 40.992 ;
 RECT 3.584 40.6035 3.64 40.8035 ;
 RECT 4.172 40.6895 4.228 40.8895 ;
 RECT 4.76 40.768 4.816 40.968 ;
 RECT 4.928 40.646 4.984 40.846 ;
 RECT 5.096 40.792 5.152 40.992 ;
 END
 END vccd_1p0.gds1669
 PIN vccd_1p0.gds1670
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 42.9965 6.838 43.1965 ;
 END
 END vccd_1p0.gds1670
 PIN vccd_1p0.gds1671
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 42.9985 5.602 43.1985 ;
 END
 END vccd_1p0.gds1671
 PIN vccd_1p0.gds1672
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 40.486 6.05 40.686 ;
 END
 END vccd_1p0.gds1672
 PIN vccd_1p0.gds1673
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 41.0165 5.41 41.2165 ;
 END
 END vccd_1p0.gds1673
 PIN vccd_1p0.gds1674
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 44.9775 5.922 45.1775 ;
 END
 END vccd_1p0.gds1674
 PIN vccd_1p0.gds1675
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.754 41.3765 5.794 41.5765 ;
 END
 END vccd_1p0.gds1675
 PIN vccd_1p0.gds1676
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 44.213 6.306 44.413 ;
 END
 END vccd_1p0.gds1676
 PIN vccd_1p0.gds1677
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 43.067 6.582 43.267 ;
 END
 END vccd_1p0.gds1677
 PIN vccd_1p0.gds1678
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.6 44.4695 5.656 44.6695 ;
 RECT 5.264 44.4695 5.32 44.6695 ;
 RECT 5.432 44.3835 5.488 44.5835 ;
 RECT 5.936 44.3835 5.992 44.5835 ;
 RECT 5.768 44.3835 5.824 44.5835 ;
 RECT 6.44 44.398 6.496 44.598 ;
 RECT 6.272 44.3835 6.328 44.5835 ;
 RECT 6.104 44.572 6.16 44.772 ;
 RECT 5.6 43.2095 5.656 43.4095 ;
 RECT 5.264 43.2095 5.32 43.4095 ;
 RECT 5.432 43.1235 5.488 43.3235 ;
 RECT 5.936 43.1235 5.992 43.3235 ;
 RECT 5.768 43.1235 5.824 43.3235 ;
 RECT 6.44 43.138 6.496 43.338 ;
 RECT 6.272 43.1235 6.328 43.3235 ;
 RECT 6.104 43.312 6.16 43.512 ;
 RECT 5.6 41.9495 5.656 42.1495 ;
 RECT 5.264 41.9495 5.32 42.1495 ;
 RECT 5.432 41.8635 5.488 42.0635 ;
 RECT 5.936 41.8635 5.992 42.0635 ;
 RECT 5.768 41.8635 5.824 42.0635 ;
 RECT 6.44 41.878 6.496 42.078 ;
 RECT 6.272 41.8635 6.328 42.0635 ;
 RECT 6.104 42.052 6.16 42.252 ;
 RECT 5.6 40.6895 5.656 40.8895 ;
 RECT 5.264 40.6895 5.32 40.8895 ;
 RECT 5.432 40.6035 5.488 40.8035 ;
 RECT 5.936 40.6035 5.992 40.8035 ;
 RECT 5.768 40.6035 5.824 40.8035 ;
 RECT 6.104 40.792 6.16 40.992 ;
 RECT 6.44 40.618 6.496 40.818 ;
 RECT 6.272 40.6035 6.328 40.8035 ;
 END
 END vccd_1p0.gds1678
 PIN vccd_1p0.gds1679
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 43.444 13.978 43.644 ;
 END
 END vccd_1p0.gds1679
 PIN vccd_1p0.gds1680
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 40.924 13.978 41.124 ;
 END
 END vccd_1p0.gds1680
 PIN vccd_1p0.gds1681
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 44.704 13.978 44.904 ;
 END
 END vccd_1p0.gds1681
 PIN vccd_1p0.gds1682
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 42.184 13.978 42.384 ;
 END
 END vccd_1p0.gds1682
 PIN vccd_1p0.gds1683
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 40.924 14.398 41.124 ;
 END
 END vccd_1p0.gds1683
 PIN vccd_1p0.gds1684
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 41.0515 14.934 41.2515 ;
 END
 END vccd_1p0.gds1684
 PIN vccd_1p0.gds1685
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 42.184 14.398 42.384 ;
 END
 END vccd_1p0.gds1685
 PIN vccd_1p0.gds1686
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 42.3115 14.934 42.5115 ;
 END
 END vccd_1p0.gds1686
 PIN vccd_1p0.gds1687
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 43.444 14.398 43.644 ;
 END
 END vccd_1p0.gds1687
 PIN vccd_1p0.gds1688
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 43.5715 14.934 43.7715 ;
 END
 END vccd_1p0.gds1688
 PIN vccd_1p0.gds1689
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 44.704 14.398 44.904 ;
 END
 END vccd_1p0.gds1689
 PIN vccd_1p0.gds1690
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 44.8315 14.934 45.0315 ;
 END
 END vccd_1p0.gds1690
 PIN vccd_1p0.gds1691
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 43.958 13.738 44.158 ;
 END
 END vccd_1p0.gds1691
 PIN vccd_1p0.gds1692
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 44.3515 13.138 44.5515 ;
 END
 END vccd_1p0.gds1692
 PIN vccd_1p0.gds1693
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 42.584 12.898 42.784 ;
 END
 END vccd_1p0.gds1693
 PIN vccd_1p0.gds1694
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 43.527 12.654 43.727 ;
 END
 END vccd_1p0.gds1694
 PIN vccd_1p0.gds1695
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 40.9985 12.526 41.1985 ;
 END
 END vccd_1p0.gds1695
 PIN vccd_1p0.gds1696
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 41.586 14.742 41.786 ;
 END
 END vccd_1p0.gds1696
 PIN vccd_1p0.gds1697
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 40.988 16.226 41.188 ;
 END
 END vccd_1p0.gds1697
 PIN vccd_1p0.gds1698
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 42.248 16.226 42.448 ;
 END
 END vccd_1p0.gds1698
 PIN vccd_1p0.gds1699
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 43.508 16.226 43.708 ;
 END
 END vccd_1p0.gds1699
 PIN vccd_1p0.gds1700
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 44.768 16.226 44.968 ;
 END
 END vccd_1p0.gds1700
 PIN vccd_1p0.gds1701
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 43.72 15.742 43.92 ;
 END
 END vccd_1p0.gds1701
 PIN vccd_1p0.gds1702
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 44.946 15.29 45.146 ;
 END
 END vccd_1p0.gds1702
 PIN vccd_1p0.gds1703
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 42.727 17.574 42.927 ;
 END
 END vccd_1p0.gds1703
 PIN vccd_1p0.gds1704
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 44.7075 18.09 44.9075 ;
 END
 END vccd_1p0.gds1704
 PIN vccd_1p0.gds1705
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 44.787 17.962 44.987 ;
 END
 END vccd_1p0.gds1705
 PIN vccd_1p0.gds1706
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 44.5235 17.734 44.7235 ;
 END
 END vccd_1p0.gds1706
 PIN vccd_1p0.gds1707
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 43.563 15.498 43.763 ;
 END
 END vccd_1p0.gds1707
 PIN vccd_1p0.gds1708
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 41.7785 17.154 41.9785 ;
 END
 END vccd_1p0.gds1708
 PIN vccd_1p0.gds1709
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 43.0675 23.842 43.2675 ;
 END
 END vccd_1p0.gds1709
 PIN vccd_1p0.gds1710
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 43.527 29.706 43.727 ;
 END
 END vccd_1p0.gds1710
 PIN vccd_1p0.gds1711
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 40.9985 29.578 41.1985 ;
 END
 END vccd_1p0.gds1711
 PIN vccd_1p0.gds1712
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 42.584 29.95 42.784 ;
 END
 END vccd_1p0.gds1712
 PIN vccd_1p0.gds1713
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 40.988 33.278 41.188 ;
 END
 END vccd_1p0.gds1713
 PIN vccd_1p0.gds1714
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 40.924 31.45 41.124 ;
 END
 END vccd_1p0.gds1714
 PIN vccd_1p0.gds1715
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 41.0515 31.986 41.2515 ;
 END
 END vccd_1p0.gds1715
 PIN vccd_1p0.gds1716
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 42.248 33.278 42.448 ;
 END
 END vccd_1p0.gds1716
 PIN vccd_1p0.gds1717
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 42.184 31.45 42.384 ;
 END
 END vccd_1p0.gds1717
 PIN vccd_1p0.gds1718
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 42.3115 31.986 42.5115 ;
 END
 END vccd_1p0.gds1718
 PIN vccd_1p0.gds1719
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 43.508 33.278 43.708 ;
 END
 END vccd_1p0.gds1719
 PIN vccd_1p0.gds1720
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 43.444 31.45 43.644 ;
 END
 END vccd_1p0.gds1720
 PIN vccd_1p0.gds1721
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 43.5715 31.986 43.7715 ;
 END
 END vccd_1p0.gds1721
 PIN vccd_1p0.gds1722
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 44.768 33.278 44.968 ;
 END
 END vccd_1p0.gds1722
 PIN vccd_1p0.gds1723
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 44.704 31.45 44.904 ;
 END
 END vccd_1p0.gds1723
 PIN vccd_1p0.gds1724
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 44.8315 31.986 45.0315 ;
 END
 END vccd_1p0.gds1724
 PIN vccd_1p0.gds1725
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 44.946 32.342 45.146 ;
 END
 END vccd_1p0.gds1725
 PIN vccd_1p0.gds1726
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 40.924 31.03 41.124 ;
 END
 END vccd_1p0.gds1726
 PIN vccd_1p0.gds1727
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 42.184 31.03 42.384 ;
 END
 END vccd_1p0.gds1727
 PIN vccd_1p0.gds1728
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 43.444 31.03 43.644 ;
 END
 END vccd_1p0.gds1728
 PIN vccd_1p0.gds1729
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 44.704 31.03 44.904 ;
 END
 END vccd_1p0.gds1729
 PIN vccd_1p0.gds1730
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 43.958 30.79 44.158 ;
 END
 END vccd_1p0.gds1730
 PIN vccd_1p0.gds1731
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 44.3515 30.19 44.5515 ;
 END
 END vccd_1p0.gds1731
 PIN vccd_1p0.gds1732
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 41.586 31.794 41.786 ;
 END
 END vccd_1p0.gds1732
 PIN vccd_1p0.gds1733
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 42.727 34.626 42.927 ;
 END
 END vccd_1p0.gds1733
 PIN vccd_1p0.gds1734
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 44.7075 35.142 44.9075 ;
 END
 END vccd_1p0.gds1734
 PIN vccd_1p0.gds1735
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 44.787 35.014 44.987 ;
 END
 END vccd_1p0.gds1735
 PIN vccd_1p0.gds1736
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 41.7785 34.206 41.9785 ;
 END
 END vccd_1p0.gds1736
 PIN vccd_1p0.gds1737
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 43.563 32.55 43.763 ;
 END
 END vccd_1p0.gds1737
 PIN vccd_1p0.gds1738
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 44.5235 34.786 44.7235 ;
 END
 END vccd_1p0.gds1738
 PIN vccd_1p0.gds1739
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 43.72 32.794 43.92 ;
 END
 END vccd_1p0.gds1739
 PIN vccd_1p0.gds1740
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 43.0675 40.894 43.2675 ;
 END
 END vccd_1p0.gds1740
 PIN vccd_1p0.gds1741
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 40.924 48.082 41.124 ;
 END
 END vccd_1p0.gds1741
 PIN vccd_1p0.gds1742
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 42.184 48.082 42.384 ;
 END
 END vccd_1p0.gds1742
 PIN vccd_1p0.gds1743
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 43.444 48.082 43.644 ;
 END
 END vccd_1p0.gds1743
 PIN vccd_1p0.gds1744
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 44.704 48.082 44.904 ;
 END
 END vccd_1p0.gds1744
 PIN vccd_1p0.gds1745
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 40.924 48.502 41.124 ;
 END
 END vccd_1p0.gds1745
 PIN vccd_1p0.gds1746
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 41.0515 49.038 41.2515 ;
 END
 END vccd_1p0.gds1746
 PIN vccd_1p0.gds1747
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 42.184 48.502 42.384 ;
 END
 END vccd_1p0.gds1747
 PIN vccd_1p0.gds1748
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 42.3115 49.038 42.5115 ;
 END
 END vccd_1p0.gds1748
 PIN vccd_1p0.gds1749
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 43.444 48.502 43.644 ;
 END
 END vccd_1p0.gds1749
 PIN vccd_1p0.gds1750
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 43.5715 49.038 43.7715 ;
 END
 END vccd_1p0.gds1750
 PIN vccd_1p0.gds1751
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 44.704 48.502 44.904 ;
 END
 END vccd_1p0.gds1751
 PIN vccd_1p0.gds1752
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 44.8315 49.038 45.0315 ;
 END
 END vccd_1p0.gds1752
 PIN vccd_1p0.gds1753
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 44.946 49.394 45.146 ;
 END
 END vccd_1p0.gds1753
 PIN vccd_1p0.gds1754
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 43.958 47.842 44.158 ;
 END
 END vccd_1p0.gds1754
 PIN vccd_1p0.gds1755
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 44.3515 47.242 44.5515 ;
 END
 END vccd_1p0.gds1755
 PIN vccd_1p0.gds1756
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 43.527 46.758 43.727 ;
 END
 END vccd_1p0.gds1756
 PIN vccd_1p0.gds1757
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 40.9985 46.63 41.1985 ;
 END
 END vccd_1p0.gds1757
 PIN vccd_1p0.gds1758
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 42.584 47.002 42.784 ;
 END
 END vccd_1p0.gds1758
 PIN vccd_1p0.gds1759
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 41.586 48.846 41.786 ;
 END
 END vccd_1p0.gds1759
 PIN vccd_1p0.gds1760
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 43.563 49.602 43.763 ;
 END
 END vccd_1p0.gds1760
 PIN vccd_1p0.gds1761
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 43.72 49.846 43.92 ;
 END
 END vccd_1p0.gds1761
 PIN vccd_1p0.gds1762
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 40.988 50.33 41.188 ;
 END
 END vccd_1p0.gds1762
 PIN vccd_1p0.gds1763
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 42.248 50.33 42.448 ;
 END
 END vccd_1p0.gds1763
 PIN vccd_1p0.gds1764
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 43.508 50.33 43.708 ;
 END
 END vccd_1p0.gds1764
 PIN vccd_1p0.gds1765
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 44.768 50.33 44.968 ;
 END
 END vccd_1p0.gds1765
 PIN vccd_1p0.gds1766
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 42.727 51.678 42.927 ;
 END
 END vccd_1p0.gds1766
 PIN vccd_1p0.gds1767
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 44.7075 52.194 44.9075 ;
 END
 END vccd_1p0.gds1767
 PIN vccd_1p0.gds1768
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 44.787 52.066 44.987 ;
 END
 END vccd_1p0.gds1768
 PIN vccd_1p0.gds1769
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 41.7785 51.258 41.9785 ;
 END
 END vccd_1p0.gds1769
 PIN vccd_1p0.gds1770
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 44.5235 51.838 44.7235 ;
 END
 END vccd_1p0.gds1770
 PIN vccd_1p0.gds1771
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 43.0675 57.946 43.2675 ;
 END
 END vccd_1p0.gds1771
 PIN vccd_1p0.gds1772
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 40.924 65.134 41.124 ;
 END
 END vccd_1p0.gds1772
 PIN vccd_1p0.gds1773
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 42.184 65.134 42.384 ;
 END
 END vccd_1p0.gds1773
 PIN vccd_1p0.gds1774
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 43.444 65.134 43.644 ;
 END
 END vccd_1p0.gds1774
 PIN vccd_1p0.gds1775
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 44.704 65.134 44.904 ;
 END
 END vccd_1p0.gds1775
 PIN vccd_1p0.gds1776
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 43.958 64.894 44.158 ;
 END
 END vccd_1p0.gds1776
 PIN vccd_1p0.gds1777
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 44.3515 64.294 44.5515 ;
 END
 END vccd_1p0.gds1777
 PIN vccd_1p0.gds1778
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 43.527 63.81 43.727 ;
 END
 END vccd_1p0.gds1778
 PIN vccd_1p0.gds1779
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 40.9985 63.682 41.1985 ;
 END
 END vccd_1p0.gds1779
 PIN vccd_1p0.gds1780
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 42.584 64.054 42.784 ;
 END
 END vccd_1p0.gds1780
 PIN vccd_1p0.gds1781
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 40.988 67.382 41.188 ;
 END
 END vccd_1p0.gds1781
 PIN vccd_1p0.gds1782
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 40.924 65.554 41.124 ;
 END
 END vccd_1p0.gds1782
 PIN vccd_1p0.gds1783
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 41.0515 66.09 41.2515 ;
 END
 END vccd_1p0.gds1783
 PIN vccd_1p0.gds1784
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 42.248 67.382 42.448 ;
 END
 END vccd_1p0.gds1784
 PIN vccd_1p0.gds1785
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 42.184 65.554 42.384 ;
 END
 END vccd_1p0.gds1785
 PIN vccd_1p0.gds1786
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 42.3115 66.09 42.5115 ;
 END
 END vccd_1p0.gds1786
 PIN vccd_1p0.gds1787
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 43.508 67.382 43.708 ;
 END
 END vccd_1p0.gds1787
 PIN vccd_1p0.gds1788
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 43.444 65.554 43.644 ;
 END
 END vccd_1p0.gds1788
 PIN vccd_1p0.gds1789
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 43.5715 66.09 43.7715 ;
 END
 END vccd_1p0.gds1789
 PIN vccd_1p0.gds1790
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 44.768 67.382 44.968 ;
 END
 END vccd_1p0.gds1790
 PIN vccd_1p0.gds1791
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 44.704 65.554 44.904 ;
 END
 END vccd_1p0.gds1791
 PIN vccd_1p0.gds1792
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 44.8315 66.09 45.0315 ;
 END
 END vccd_1p0.gds1792
 PIN vccd_1p0.gds1793
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 44.946 66.446 45.146 ;
 END
 END vccd_1p0.gds1793
 PIN vccd_1p0.gds1794
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 41.586 65.898 41.786 ;
 END
 END vccd_1p0.gds1794
 PIN vccd_1p0.gds1795
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 42.727 68.73 42.927 ;
 END
 END vccd_1p0.gds1795
 PIN vccd_1p0.gds1796
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 44.7075 69.246 44.9075 ;
 END
 END vccd_1p0.gds1796
 PIN vccd_1p0.gds1797
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 44.787 69.118 44.987 ;
 END
 END vccd_1p0.gds1797
 PIN vccd_1p0.gds1798
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 41.7785 68.31 41.9785 ;
 END
 END vccd_1p0.gds1798
 PIN vccd_1p0.gds1799
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 43.563 66.654 43.763 ;
 END
 END vccd_1p0.gds1799
 PIN vccd_1p0.gds1800
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 44.5235 68.89 44.7235 ;
 END
 END vccd_1p0.gds1800
 PIN vccd_1p0.gds1801
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 43.72 66.898 43.92 ;
 END
 END vccd_1p0.gds1801
 PIN vccd_1p0.gds1802
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.384 47.199 0.43 47.399 ;
 END
 END vccd_1p0.gds1802
 PIN vccd_1p0.gds1803
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 46.0245 4.738 46.2245 ;
 END
 END vccd_1p0.gds1803
 PIN vccd_1p0.gds1804
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.698 48.687 4.738 48.887 ;
 END
 END vccd_1p0.gds1804
 PIN vccd_1p0.gds1805
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 48.137 1.542 48.337 ;
 END
 END vccd_1p0.gds1805
 PIN vccd_1p0.gds1806
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 48.109 5.202 48.309 ;
 END
 END vccd_1p0.gds1806
 PIN vccd_1p0.gds1807
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 46.877 1.542 47.077 ;
 END
 END vccd_1p0.gds1807
 PIN vccd_1p0.gds1808
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.486 45.617 1.542 45.817 ;
 END
 END vccd_1p0.gds1808
 PIN vccd_1p0.gds1809
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.518 47.36 0.548 47.56 ;
 END
 END vccd_1p0.gds1809
 PIN vccd_1p0.gds1810
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.726 47.968 1.782 48.168 ;
 END
 END vccd_1p0.gds1810
 PIN vccd_1p0.gds1811
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 0.812 47.183 0.858 47.383 ;
 END
 END vccd_1p0.gds1811
 PIN vccd_1p0.gds1812
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.306 47.314 1.362 47.514 ;
 END
 END vccd_1p0.gds1812
 PIN vccd_1p0.gds1813
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.178 47.2975 1.218 47.4975 ;
 END
 END vccd_1p0.gds1813
 PIN vccd_1p0.gds1814
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.05 47.211 1.09 47.411 ;
 END
 END vccd_1p0.gds1814
 PIN vccd_1p0.gds1815
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.146 48.328 2.202 48.528 ;
 END
 END vccd_1p0.gds1815
 PIN vccd_1p0.gds1816
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.566 47.152 2.622 47.352 ;
 END
 END vccd_1p0.gds1816
 PIN vccd_1p0.gds1817
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.406 48.377 2.462 48.577 ;
 END
 END vccd_1p0.gds1817
 PIN vccd_1p0.gds1818
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 45.4995 5.202 45.6995 ;
 END
 END vccd_1p0.gds1818
 PIN vccd_1p0.gds1819
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.986 47.1825 3.042 47.3825 ;
 END
 END vccd_1p0.gds1819
 PIN vccd_1p0.gds1820
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.162 46.7595 5.202 46.9595 ;
 END
 END vccd_1p0.gds1820
 PIN vccd_1p0.gds1821
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 1.906 47.131 1.962 47.331 ;
 END
 END vccd_1p0.gds1821
 PIN vccd_1p0.gds1822
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 2.826 47.258 2.882 47.458 ;
 END
 END vccd_1p0.gds1822
 PIN vccd_1p0.gds1823
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.35 47.2825 3.39 47.4825 ;
 END
 END vccd_1p0.gds1823
 PIN vccd_1p0.gds1824
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.23 47.2035 3.262 47.4035 ;
 END
 END vccd_1p0.gds1824
 PIN vccd_1p0.gds1825
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 48.7075 3.666 48.9075 ;
 END
 END vccd_1p0.gds1825
 PIN vccd_1p0.gds1826
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.626 45.983 3.666 46.183 ;
 END
 END vccd_1p0.gds1826
 PIN vccd_1p0.gds1827
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 48.58 4.066 48.78 ;
 END
 END vccd_1p0.gds1827
 PIN vccd_1p0.gds1828
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.026 45.6965 4.066 45.8965 ;
 END
 END vccd_1p0.gds1828
 PIN vccd_1p0.gds1829
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.218 46.6245 4.258 46.8245 ;
 END
 END vccd_1p0.gds1829
 PIN vccd_1p0.gds1830
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 3.818 47.2325 3.858 47.4325 ;
 END
 END vccd_1p0.gds1830
 PIN vccd_1p0.gds1831
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.506 47.2415 4.546 47.4415 ;
 END
 END vccd_1p0.gds1831
 PIN vccd_1p0.gds1832
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 4.97 47.2395 5.01 47.4395 ;
 END
 END vccd_1p0.gds1832
 PIN vccd_1p0.gds1833
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 4.34 45.832 4.396 46.032 ;
 RECT 4.76 45.808 4.816 46.008 ;
 RECT 5.096 45.832 5.152 46.032 ;
 RECT 4.34 47.092 4.396 47.292 ;
 RECT 4.76 47.068 4.816 47.268 ;
 RECT 5.096 47.092 5.152 47.292 ;
 RECT 4.34 48.352 4.396 48.552 ;
 RECT 4.76 48.328 4.816 48.528 ;
 RECT 5.096 48.352 5.152 48.552 ;
 RECT 3.584 48.1635 3.64 48.3635 ;
 RECT 4.172 48.2495 4.228 48.4495 ;
 RECT 4.928 48.206 4.984 48.406 ;
 RECT 3.584 46.9035 3.64 47.1035 ;
 RECT 4.172 46.9895 4.228 47.1895 ;
 RECT 4.928 46.946 4.984 47.146 ;
 RECT 3.584 45.6435 3.64 45.8435 ;
 RECT 4.172 45.7295 4.228 45.9295 ;
 RECT 4.928 45.686 4.984 45.886 ;
 END
 END vccd_1p0.gds1833
 PIN vccd_1p0.gds1834
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.798 47.2325 6.838 47.4325 ;
 END
 END vccd_1p0.gds1834
 PIN vccd_1p0.gds1835
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.562 47.171 5.602 47.371 ;
 END
 END vccd_1p0.gds1835
 PIN vccd_1p0.gds1836
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 48.5095 6.05 48.7095 ;
 END
 END vccd_1p0.gds1836
 PIN vccd_1p0.gds1837
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.01 45.526 6.05 45.726 ;
 END
 END vccd_1p0.gds1837
 PIN vccd_1p0.gds1838
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 48.644 5.41 48.844 ;
 END
 END vccd_1p0.gds1838
 PIN vccd_1p0.gds1839
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.37 45.965 5.41 46.165 ;
 END
 END vccd_1p0.gds1839
 PIN vccd_1p0.gds1840
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.882 48.13 5.922 48.33 ;
 END
 END vccd_1p0.gds1840
 PIN vccd_1p0.gds1841
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 5.754 46.4165 5.794 46.6165 ;
 END
 END vccd_1p0.gds1841
 PIN vccd_1p0.gds1842
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.266 47.856 6.306 48.056 ;
 END
 END vccd_1p0.gds1842
 PIN vccd_1p0.gds1843
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 6.522 47.2285 6.582 47.4285 ;
 END
 END vccd_1p0.gds1843
 PIN vccd_1p0.gds1844
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 5.6 48.2495 5.656 48.4495 ;
 RECT 5.264 48.2495 5.32 48.4495 ;
 RECT 5.432 48.1635 5.488 48.3635 ;
 RECT 5.936 48.1635 5.992 48.3635 ;
 RECT 5.768 48.1635 5.824 48.3635 ;
 RECT 6.44 48.178 6.496 48.378 ;
 RECT 6.272 48.1635 6.328 48.3635 ;
 RECT 6.104 48.352 6.16 48.552 ;
 RECT 5.6 46.9895 5.656 47.1895 ;
 RECT 5.264 46.9895 5.32 47.1895 ;
 RECT 5.432 46.9035 5.488 47.1035 ;
 RECT 5.936 46.9035 5.992 47.1035 ;
 RECT 5.768 46.9035 5.824 47.1035 ;
 RECT 6.44 46.918 6.496 47.118 ;
 RECT 6.272 46.9035 6.328 47.1035 ;
 RECT 6.104 47.092 6.16 47.292 ;
 RECT 5.6 45.7295 5.656 45.9295 ;
 RECT 5.264 45.7295 5.32 45.9295 ;
 RECT 5.432 45.6435 5.488 45.8435 ;
 RECT 5.936 45.6435 5.992 45.8435 ;
 RECT 5.768 45.6435 5.824 45.8435 ;
 RECT 6.44 45.658 6.496 45.858 ;
 RECT 6.272 45.6435 6.328 45.8435 ;
 RECT 6.104 45.832 6.16 46.032 ;
 END
 END vccd_1p0.gds1844
 PIN vccd_1p0.gds1845
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 45.964 13.978 46.164 ;
 END
 END vccd_1p0.gds1845
 PIN vccd_1p0.gds1846
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 47.224 13.978 47.424 ;
 END
 END vccd_1p0.gds1846
 PIN vccd_1p0.gds1847
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.922 48.484 13.978 48.684 ;
 END
 END vccd_1p0.gds1847
 PIN vccd_1p0.gds1848
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 47.224 14.398 47.424 ;
 END
 END vccd_1p0.gds1848
 PIN vccd_1p0.gds1849
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.682 47.5135 13.738 47.7135 ;
 END
 END vccd_1p0.gds1849
 PIN vccd_1p0.gds1850
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 13.082 47.8075 13.138 48.0075 ;
 END
 END vccd_1p0.gds1850
 PIN vccd_1p0.gds1851
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.842 46.994 12.898 47.194 ;
 END
 END vccd_1p0.gds1851
 PIN vccd_1p0.gds1852
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.614 47.406 12.654 47.606 ;
 END
 END vccd_1p0.gds1852
 PIN vccd_1p0.gds1853
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 48.7075 12.526 48.9075 ;
 END
 END vccd_1p0.gds1853
 PIN vccd_1p0.gds1854
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 12.486 46.0385 12.526 46.2385 ;
 END
 END vccd_1p0.gds1854
 PIN vccd_1p0.gds1855
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 45.964 14.398 46.164 ;
 END
 END vccd_1p0.gds1855
 PIN vccd_1p0.gds1856
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 46.0915 14.934 46.2915 ;
 END
 END vccd_1p0.gds1856
 PIN vccd_1p0.gds1857
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.342 48.484 14.398 48.684 ;
 END
 END vccd_1p0.gds1857
 PIN vccd_1p0.gds1858
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 48.6115 14.934 48.8115 ;
 END
 END vccd_1p0.gds1858
 PIN vccd_1p0.gds1859
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.682 46.524 14.742 46.724 ;
 END
 END vccd_1p0.gds1859
 PIN vccd_1p0.gds1860
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 14.894 47.3515 14.934 47.5515 ;
 END
 END vccd_1p0.gds1860
 PIN vccd_1p0.gds1861
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 47.288 16.226 47.488 ;
 END
 END vccd_1p0.gds1861
 PIN vccd_1p0.gds1862
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 48.548 16.226 48.748 ;
 END
 END vccd_1p0.gds1862
 PIN vccd_1p0.gds1863
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 16.17 46.028 16.226 46.228 ;
 END
 END vccd_1p0.gds1863
 PIN vccd_1p0.gds1864
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.686 47.5015 15.742 47.7015 ;
 END
 END vccd_1p0.gds1864
 PIN vccd_1p0.gds1865
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.25 48.192 15.29 48.392 ;
 END
 END vccd_1p0.gds1865
 PIN vccd_1p0.gds1866
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.518 46.994 17.574 47.194 ;
 END
 END vccd_1p0.gds1866
 PIN vccd_1p0.gds1867
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 18.05 48.0025 18.09 48.2025 ;
 END
 END vccd_1p0.gds1867
 PIN vccd_1p0.gds1868
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.922 48.033 17.962 48.233 ;
 END
 END vccd_1p0.gds1868
 PIN vccd_1p0.gds1869
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.678 47.9475 17.734 48.1475 ;
 END
 END vccd_1p0.gds1869
 PIN vccd_1p0.gds1870
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 15.442 47.5015 15.498 47.7015 ;
 END
 END vccd_1p0.gds1870
 PIN vccd_1p0.gds1871
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 17.098 46.536 17.154 46.736 ;
 END
 END vccd_1p0.gds1871
 PIN vccd_1p0.gds1872
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 23.786 47.219 23.842 47.419 ;
 END
 END vccd_1p0.gds1872
 PIN vccd_1p0.gds1873
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.666 47.406 29.706 47.606 ;
 END
 END vccd_1p0.gds1873
 PIN vccd_1p0.gds1874
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 48.7075 29.578 48.9075 ;
 END
 END vccd_1p0.gds1874
 PIN vccd_1p0.gds1875
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.538 46.0385 29.578 46.2385 ;
 END
 END vccd_1p0.gds1875
 PIN vccd_1p0.gds1876
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 29.894 46.994 29.95 47.194 ;
 END
 END vccd_1p0.gds1876
 PIN vccd_1p0.gds1877
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 47.224 31.03 47.424 ;
 END
 END vccd_1p0.gds1877
 PIN vccd_1p0.gds1878
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 47.288 33.278 47.488 ;
 END
 END vccd_1p0.gds1878
 PIN vccd_1p0.gds1879
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 47.224 31.45 47.424 ;
 END
 END vccd_1p0.gds1879
 PIN vccd_1p0.gds1880
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 48.548 33.278 48.748 ;
 END
 END vccd_1p0.gds1880
 PIN vccd_1p0.gds1881
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 48.484 31.03 48.684 ;
 END
 END vccd_1p0.gds1881
 PIN vccd_1p0.gds1882
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.974 45.964 31.03 46.164 ;
 END
 END vccd_1p0.gds1882
 PIN vccd_1p0.gds1883
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 33.222 46.028 33.278 46.228 ;
 END
 END vccd_1p0.gds1883
 PIN vccd_1p0.gds1884
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 45.964 31.45 46.164 ;
 END
 END vccd_1p0.gds1884
 PIN vccd_1p0.gds1885
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 46.0915 31.986 46.2915 ;
 END
 END vccd_1p0.gds1885
 PIN vccd_1p0.gds1886
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.302 48.192 32.342 48.392 ;
 END
 END vccd_1p0.gds1886
 PIN vccd_1p0.gds1887
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.734 47.5135 30.79 47.7135 ;
 END
 END vccd_1p0.gds1887
 PIN vccd_1p0.gds1888
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 30.134 47.8075 30.19 48.0075 ;
 END
 END vccd_1p0.gds1888
 PIN vccd_1p0.gds1889
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.734 46.524 31.794 46.724 ;
 END
 END vccd_1p0.gds1889
 PIN vccd_1p0.gds1890
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.394 48.484 31.45 48.684 ;
 END
 END vccd_1p0.gds1890
 PIN vccd_1p0.gds1891
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 48.6115 31.986 48.8115 ;
 END
 END vccd_1p0.gds1891
 PIN vccd_1p0.gds1892
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.57 46.994 34.626 47.194 ;
 END
 END vccd_1p0.gds1892
 PIN vccd_1p0.gds1893
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 35.102 48.0025 35.142 48.2025 ;
 END
 END vccd_1p0.gds1893
 PIN vccd_1p0.gds1894
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.974 48.033 35.014 48.233 ;
 END
 END vccd_1p0.gds1894
 PIN vccd_1p0.gds1895
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.15 46.536 34.206 46.736 ;
 END
 END vccd_1p0.gds1895
 PIN vccd_1p0.gds1896
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 31.946 47.3515 31.986 47.5515 ;
 END
 END vccd_1p0.gds1896
 PIN vccd_1p0.gds1897
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.494 47.5015 32.55 47.7015 ;
 END
 END vccd_1p0.gds1897
 PIN vccd_1p0.gds1898
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 34.73 47.9475 34.786 48.1475 ;
 END
 END vccd_1p0.gds1898
 PIN vccd_1p0.gds1899
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 32.738 47.5015 32.794 47.7015 ;
 END
 END vccd_1p0.gds1899
 PIN vccd_1p0.gds1900
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 40.838 47.219 40.894 47.419 ;
 END
 END vccd_1p0.gds1900
 PIN vccd_1p0.gds1901
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 47.224 48.082 47.424 ;
 END
 END vccd_1p0.gds1901
 PIN vccd_1p0.gds1902
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 48.484 48.082 48.684 ;
 END
 END vccd_1p0.gds1902
 PIN vccd_1p0.gds1903
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 47.224 48.502 47.424 ;
 END
 END vccd_1p0.gds1903
 PIN vccd_1p0.gds1904
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.026 45.964 48.082 46.164 ;
 END
 END vccd_1p0.gds1904
 PIN vccd_1p0.gds1905
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 45.964 48.502 46.164 ;
 END
 END vccd_1p0.gds1905
 PIN vccd_1p0.gds1906
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 46.0915 49.038 46.2915 ;
 END
 END vccd_1p0.gds1906
 PIN vccd_1p0.gds1907
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.354 48.192 49.394 48.392 ;
 END
 END vccd_1p0.gds1907
 PIN vccd_1p0.gds1908
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.786 47.5135 47.842 47.7135 ;
 END
 END vccd_1p0.gds1908
 PIN vccd_1p0.gds1909
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 47.186 47.8075 47.242 48.0075 ;
 END
 END vccd_1p0.gds1909
 PIN vccd_1p0.gds1910
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.718 47.406 46.758 47.606 ;
 END
 END vccd_1p0.gds1910
 PIN vccd_1p0.gds1911
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 48.7075 46.63 48.9075 ;
 END
 END vccd_1p0.gds1911
 PIN vccd_1p0.gds1912
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.59 46.0385 46.63 46.2385 ;
 END
 END vccd_1p0.gds1912
 PIN vccd_1p0.gds1913
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 46.946 46.994 47.002 47.194 ;
 END
 END vccd_1p0.gds1913
 PIN vccd_1p0.gds1914
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.786 46.524 48.846 46.724 ;
 END
 END vccd_1p0.gds1914
 PIN vccd_1p0.gds1915
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.446 48.484 48.502 48.684 ;
 END
 END vccd_1p0.gds1915
 PIN vccd_1p0.gds1916
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 48.6115 49.038 48.8115 ;
 END
 END vccd_1p0.gds1916
 PIN vccd_1p0.gds1917
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 48.998 47.3515 49.038 47.5515 ;
 END
 END vccd_1p0.gds1917
 PIN vccd_1p0.gds1918
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.546 47.5015 49.602 47.7015 ;
 END
 END vccd_1p0.gds1918
 PIN vccd_1p0.gds1919
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 49.79 47.5015 49.846 47.7015 ;
 END
 END vccd_1p0.gds1919
 PIN vccd_1p0.gds1920
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 47.288 50.33 47.488 ;
 END
 END vccd_1p0.gds1920
 PIN vccd_1p0.gds1921
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 48.548 50.33 48.748 ;
 END
 END vccd_1p0.gds1921
 PIN vccd_1p0.gds1922
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 50.274 46.028 50.33 46.228 ;
 END
 END vccd_1p0.gds1922
 PIN vccd_1p0.gds1923
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.622 46.994 51.678 47.194 ;
 END
 END vccd_1p0.gds1923
 PIN vccd_1p0.gds1924
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.154 48.0025 52.194 48.2025 ;
 END
 END vccd_1p0.gds1924
 PIN vccd_1p0.gds1925
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 52.026 48.033 52.066 48.233 ;
 END
 END vccd_1p0.gds1925
 PIN vccd_1p0.gds1926
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.202 46.536 51.258 46.736 ;
 END
 END vccd_1p0.gds1926
 PIN vccd_1p0.gds1927
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 51.782 47.9475 51.838 48.1475 ;
 END
 END vccd_1p0.gds1927
 PIN vccd_1p0.gds1928
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 57.89 47.219 57.946 47.419 ;
 END
 END vccd_1p0.gds1928
 PIN vccd_1p0.gds1929
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 47.224 65.134 47.424 ;
 END
 END vccd_1p0.gds1929
 PIN vccd_1p0.gds1930
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 48.484 65.134 48.684 ;
 END
 END vccd_1p0.gds1930
 PIN vccd_1p0.gds1931
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.078 45.964 65.134 46.164 ;
 END
 END vccd_1p0.gds1931
 PIN vccd_1p0.gds1932
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.838 47.5135 64.894 47.7135 ;
 END
 END vccd_1p0.gds1932
 PIN vccd_1p0.gds1933
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 64.238 47.8075 64.294 48.0075 ;
 END
 END vccd_1p0.gds1933
 PIN vccd_1p0.gds1934
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.77 47.406 63.81 47.606 ;
 END
 END vccd_1p0.gds1934
 PIN vccd_1p0.gds1935
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 48.7075 63.682 48.9075 ;
 END
 END vccd_1p0.gds1935
 PIN vccd_1p0.gds1936
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.642 46.0385 63.682 46.2385 ;
 END
 END vccd_1p0.gds1936
 PIN vccd_1p0.gds1937
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 63.998 46.994 64.054 47.194 ;
 END
 END vccd_1p0.gds1937
 PIN vccd_1p0.gds1938
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 47.288 67.382 47.488 ;
 END
 END vccd_1p0.gds1938
 PIN vccd_1p0.gds1939
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 47.224 65.554 47.424 ;
 END
 END vccd_1p0.gds1939
 PIN vccd_1p0.gds1940
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 48.548 67.382 48.748 ;
 END
 END vccd_1p0.gds1940
 PIN vccd_1p0.gds1941
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 67.326 46.028 67.382 46.228 ;
 END
 END vccd_1p0.gds1941
 PIN vccd_1p0.gds1942
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 45.964 65.554 46.164 ;
 END
 END vccd_1p0.gds1942
 PIN vccd_1p0.gds1943
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 46.0915 66.09 46.2915 ;
 END
 END vccd_1p0.gds1943
 PIN vccd_1p0.gds1944
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.406 48.192 66.446 48.392 ;
 END
 END vccd_1p0.gds1944
 PIN vccd_1p0.gds1945
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.838 46.524 65.898 46.724 ;
 END
 END vccd_1p0.gds1945
 PIN vccd_1p0.gds1946
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 65.498 48.484 65.554 48.684 ;
 END
 END vccd_1p0.gds1946
 PIN vccd_1p0.gds1947
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 48.6115 66.09 48.8115 ;
 END
 END vccd_1p0.gds1947
 PIN vccd_1p0.gds1948
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.674 46.994 68.73 47.194 ;
 END
 END vccd_1p0.gds1948
 PIN vccd_1p0.gds1949
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.206 48.0025 69.246 48.2025 ;
 END
 END vccd_1p0.gds1949
 PIN vccd_1p0.gds1950
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 69.078 48.033 69.118 48.233 ;
 END
 END vccd_1p0.gds1950
 PIN vccd_1p0.gds1951
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.254 46.536 68.31 46.736 ;
 END
 END vccd_1p0.gds1951
 PIN vccd_1p0.gds1952
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.05 47.3515 66.09 47.5515 ;
 END
 END vccd_1p0.gds1952
 PIN vccd_1p0.gds1953
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.598 47.5015 66.654 47.7015 ;
 END
 END vccd_1p0.gds1953
 PIN vccd_1p0.gds1954
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 68.834 47.9475 68.89 48.1475 ;
 END
 END vccd_1p0.gds1954
 PIN vccd_1p0.gds1955
 DIRECTION INPUT ;
 USE POWER ;
 PORT
 LAYER m3 ;
 RECT 66.842 47.5015 66.898 47.7015 ;
 END
 END vccd_1p0.gds1955
 PIN vss
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 0.913 2.962 1.113 ;
 END
 END vss
 PIN vss.gds1
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 2.173 2.962 2.373 ;
 END
 END vss.gds1
 PIN vss.gds2
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 3.433 2.962 3.633 ;
 END
 END vss.gds2
 PIN vss.gds3
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 0.6075 3.142 0.8075 ;
 END
 END vss.gds3
 PIN vss.gds4
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 4.693 2.962 4.893 ;
 END
 END vss.gds4
 PIN vss.gds5
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 2.397 0.942 2.597 ;
 END
 END vss.gds5
 PIN vss.gds6
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.286 2.803 3.326 3.003 ;
 END
 END vss.gds6
 PIN vss.gds7
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 2.803 4.194 3.003 ;
 END
 END vss.gds7
 PIN vss.gds8
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 2.803 5.074 3.003 ;
 END
 END vss.gds8
 PIN vss.gds9
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 4.292 3.142 4.492 ;
 END
 END vss.gds9
 PIN vss.gds10
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 3.032 3.142 3.232 ;
 END
 END vss.gds10
 PIN vss.gds11
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 2.4975 0.718 2.6975 ;
 END
 END vss.gds11
 PIN vss.gds12
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.442 2.397 4.482 2.597 ;
 END
 END vss.gds12
 PIN vss.gds13
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.57 2.6 4.61 2.8 ;
 END
 END vss.gds13
 PIN vss.gds14
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 2.397 4.882 2.597 ;
 END
 END vss.gds14
 PIN vss.gds15
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 2.598 0.602 2.798 ;
 END
 END vss.gds15
 PIN vss.gds16
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 1.772 3.142 1.972 ;
 END
 END vss.gds16
 PIN vss.gds17
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 2.8265 2.122 3.0265 ;
 END
 END vss.gds17
 PIN vss.gds18
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 2.941 1.282 3.141 ;
 END
 END vss.gds18
 PIN vss.gds19
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 3.1755 1.462 3.3755 ;
 END
 END vss.gds19
 PIN vss.gds20
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.414 3.079 3.454 3.279 ;
 END
 END vss.gds20
 PIN vss.gds21
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.562 3.079 3.602 3.279 ;
 END
 END vss.gds21
 PIN vss.gds22
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 2.738 2.302 2.938 ;
 END
 END vss.gds22
 PIN vss.gds23
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 2.6995 4.002 2.8995 ;
 END
 END vss.gds23
 PIN vss.gds24
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 2.6995 5.282 2.8995 ;
 END
 END vss.gds24
 PIN vss.gds25
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 2.476 0.29 2.676 ;
 END
 END vss.gds25
 PIN vss.gds26
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.754 2.803 3.794 3.003 ;
 END
 END vss.gds26
 PIN vss.gds27
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 2.576 2.1735 2.632 2.3735 ;
 RECT 2.408 2.1735 2.464 2.3735 ;
 RECT 2.996 2.1735 3.052 2.3735 ;
 RECT 3.332 2.265 3.388 2.465 ;
 RECT 2.408 0.9135 2.464 1.1135 ;
 RECT 2.576 0.9135 2.632 1.1135 ;
 RECT 2.996 0.9135 3.052 1.1135 ;
 RECT 3.332 1.005 3.388 1.205 ;
 RECT 3.5 0.9615 3.556 1.1615 ;
 RECT 0.98 0.8285 1.036 1.0285 ;
 RECT 2.072 0.829 2.128 1.029 ;
 RECT 0.812 2.265 0.868 2.465 ;
 RECT 2.408 3.4335 2.464 3.6335 ;
 RECT 2.576 3.4335 2.632 3.6335 ;
 RECT 2.996 3.4335 3.052 3.6335 ;
 RECT 3.332 3.525 3.388 3.725 ;
 RECT 3.5 3.4815 3.556 3.6815 ;
 RECT 0.98 3.3485 1.036 3.5485 ;
 RECT 2.072 3.349 2.128 3.549 ;
 RECT 2.408 4.6935 2.464 4.8935 ;
 RECT 2.576 4.6935 2.632 4.8935 ;
 RECT 2.996 4.6935 3.052 4.8935 ;
 RECT 0.812 4.785 0.868 4.985 ;
 RECT 3.332 4.785 3.388 4.985 ;
 RECT 3.5 4.7415 3.556 4.9415 ;
 RECT 0.392 4.699 0.448 4.899 ;
 RECT 0.644 4.699 0.7 4.899 ;
 RECT 1.232 4.699 1.288 4.899 ;
 RECT 0.98 4.6085 1.036 4.8085 ;
 RECT 1.4 4.699 1.456 4.899 ;
 RECT 1.568 4.699 1.624 4.899 ;
 RECT 2.072 4.609 2.128 4.809 ;
 RECT 1.82 4.699 1.876 4.899 ;
 RECT 2.744 4.609 2.8 4.809 ;
 RECT 3.164 4.699 3.22 4.899 ;
 RECT 3.92 4.699 3.976 4.899 ;
 RECT 3.752 4.969 3.808 5.169 ;
 RECT 4.508 4.8985 4.564 5.0985 ;
 RECT 2.24 4.699 2.296 4.899 ;
 RECT 0.392 3.439 0.448 3.639 ;
 RECT 0.812 3.525 0.868 3.725 ;
 RECT 0.644 3.439 0.7 3.639 ;
 RECT 1.232 3.439 1.288 3.639 ;
 RECT 1.4 3.439 1.456 3.639 ;
 RECT 1.568 3.439 1.624 3.639 ;
 RECT 1.82 3.439 1.876 3.639 ;
 RECT 2.24 3.439 2.296 3.639 ;
 RECT 2.744 3.349 2.8 3.549 ;
 RECT 3.164 3.439 3.22 3.639 ;
 RECT 3.92 3.439 3.976 3.639 ;
 RECT 3.752 3.709 3.808 3.909 ;
 RECT 4.508 3.6385 4.564 3.8385 ;
 RECT 3.5 2.2215 3.556 2.4215 ;
 RECT 0.392 2.179 0.448 2.379 ;
 RECT 0.644 2.179 0.7 2.379 ;
 RECT 1.232 2.179 1.288 2.379 ;
 RECT 0.98 2.0885 1.036 2.2885 ;
 RECT 1.4 2.179 1.456 2.379 ;
 RECT 1.568 2.179 1.624 2.379 ;
 RECT 2.072 2.089 2.128 2.289 ;
 RECT 1.82 2.179 1.876 2.379 ;
 RECT 2.744 2.089 2.8 2.289 ;
 RECT 3.164 2.179 3.22 2.379 ;
 RECT 2.24 2.179 2.296 2.379 ;
 RECT 0.392 0.919 0.448 1.119 ;
 RECT 0.812 1.005 0.868 1.205 ;
 RECT 0.644 0.919 0.7 1.119 ;
 RECT 1.232 0.919 1.288 1.119 ;
 RECT 1.4 0.919 1.456 1.119 ;
 RECT 1.568 0.919 1.624 1.119 ;
 RECT 1.82 0.919 1.876 1.119 ;
 RECT 2.24 0.919 2.296 1.119 ;
 RECT 2.744 0.829 2.8 1.029 ;
 RECT 3.164 0.919 3.22 1.119 ;
 RECT 3.92 0.919 3.976 1.119 ;
 RECT 3.752 1.189 3.808 1.389 ;
 RECT 4.508 1.1185 4.564 1.3185 ;
 RECT 3.92 2.179 3.976 2.379 ;
 RECT 3.752 2.449 3.808 2.649 ;
 RECT 4.508 2.3785 4.564 2.5785 ;
 END
 END vss.gds27
 PIN vss.gds28
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.134 2.9095 10.194 3.1095 ;
 END
 END vss.gds28
 PIN vss.gds29
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.966 2.9095 10.026 3.1095 ;
 END
 END vss.gds29
 PIN vss.gds30
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.798 2.9095 9.858 3.1095 ;
 END
 END vss.gds30
 PIN vss.gds31
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 2.9095 9.69 3.1095 ;
 END
 END vss.gds31
 PIN vss.gds32
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.462 2.9095 9.522 3.1095 ;
 END
 END vss.gds32
 PIN vss.gds33
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 2.9095 9.018 3.1095 ;
 END
 END vss.gds33
 PIN vss.gds34
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.79 2.9095 8.85 3.1095 ;
 END
 END vss.gds34
 PIN vss.gds35
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.622 2.9095 8.682 3.1095 ;
 END
 END vss.gds35
 PIN vss.gds36
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.454 2.9095 8.514 3.1095 ;
 END
 END vss.gds36
 PIN vss.gds37
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 2.803 5.474 3.003 ;
 END
 END vss.gds37
 PIN vss.gds38
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 2.9095 8.346 3.1095 ;
 END
 END vss.gds38
 PIN vss.gds39
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.118 2.9095 8.178 3.1095 ;
 END
 END vss.gds39
 PIN vss.gds40
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.95 2.9095 8.01 3.1095 ;
 END
 END vss.gds40
 PIN vss.gds41
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.294 2.9095 9.354 3.1095 ;
 END
 END vss.gds41
 PIN vss.gds42
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.782 2.9095 7.842 3.1095 ;
 END
 END vss.gds42
 PIN vss.gds43
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 2.9095 7.674 3.1095 ;
 END
 END vss.gds43
 PIN vss.gds44
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.126 2.9095 9.186 3.1095 ;
 END
 END vss.gds44
 PIN vss.gds45
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.446 2.9095 7.506 3.1095 ;
 END
 END vss.gds45
 PIN vss.gds46
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.278 2.9095 7.338 3.1095 ;
 END
 END vss.gds46
 PIN vss.gds47
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.11 2.9095 7.17 3.1095 ;
 END
 END vss.gds47
 PIN vss.gds48
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 2.803 5.73 3.003 ;
 END
 END vss.gds48
 PIN vss.gds49
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 2.803 5.986 3.003 ;
 END
 END vss.gds49
 PIN vss.gds50
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 2.599 6.434 2.799 ;
 END
 END vss.gds50
 PIN vss.gds51
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 2.6 6.178 2.8 ;
 END
 END vss.gds51
 PIN vss.gds52
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 6.692 4.842 6.748 5.042 ;
 RECT 6.608 4.969 6.664 5.169 ;
 RECT 6.524 4.692 6.58 4.892 ;
 RECT 6.608 3.709 6.664 3.909 ;
 RECT 6.524 3.432 6.58 3.632 ;
 RECT 6.692 3.582 6.748 3.782 ;
 RECT 6.608 1.189 6.664 1.389 ;
 RECT 6.524 0.912 6.58 1.112 ;
 RECT 6.692 1.062 6.748 1.262 ;
 RECT 6.692 2.322 6.748 2.522 ;
 RECT 6.524 2.172 6.58 2.372 ;
 RECT 6.608 2.449 6.664 2.649 ;
 END
 END vss.gds52
 PIN vss.gds53
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 1.458 14.87 1.658 ;
 END
 END vss.gds53
 PIN vss.gds54
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 5.198 13.898 5.398 ;
 END
 END vss.gds54
 PIN vss.gds55
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 5.238 14.87 5.438 ;
 END
 END vss.gds55
 PIN vss.gds56
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 2.678 13.898 2.878 ;
 END
 END vss.gds56
 PIN vss.gds57
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 2.718 14.87 2.918 ;
 END
 END vss.gds57
 PIN vss.gds58
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 3.938 13.898 4.138 ;
 END
 END vss.gds58
 PIN vss.gds59
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 3.978 14.87 4.178 ;
 END
 END vss.gds59
 PIN vss.gds60
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.15 2.9095 12.21 3.1095 ;
 END
 END vss.gds60
 PIN vss.gds61
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.982 2.9095 12.042 3.1095 ;
 END
 END vss.gds61
 PIN vss.gds62
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.814 2.9095 11.874 3.1095 ;
 END
 END vss.gds62
 PIN vss.gds63
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.478 2.9095 11.538 3.1095 ;
 END
 END vss.gds63
 PIN vss.gds64
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.31 2.9095 11.37 3.1095 ;
 END
 END vss.gds64
 PIN vss.gds65
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 3.0755 13.058 3.2755 ;
 END
 END vss.gds65
 PIN vss.gds66
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 2.9095 11.706 3.1095 ;
 END
 END vss.gds66
 PIN vss.gds67
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.142 2.9095 11.202 3.1095 ;
 END
 END vss.gds67
 PIN vss.gds68
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.806 2.9095 10.866 3.1095 ;
 END
 END vss.gds68
 PIN vss.gds69
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.638 2.9095 10.698 3.1095 ;
 END
 END vss.gds69
 PIN vss.gds70
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.47 2.9095 10.53 3.1095 ;
 END
 END vss.gds70
 PIN vss.gds71
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 2.9095 11.034 3.1095 ;
 END
 END vss.gds71
 PIN vss.gds72
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 2.9095 10.362 3.1095 ;
 END
 END vss.gds72
 PIN vss.gds73
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 3.06 15.162 3.26 ;
 END
 END vss.gds73
 PIN vss.gds74
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 3.06 14.498 3.26 ;
 END
 END vss.gds74
 PIN vss.gds75
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 3.0195 13.658 3.2195 ;
 END
 END vss.gds75
 PIN vss.gds76
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.262 3.072 13.318 3.272 ;
 END
 END vss.gds76
 PIN vss.gds77
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 2.941 12.378 3.141 ;
 END
 END vss.gds77
 PIN vss.gds78
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 2.803 12.59 3.003 ;
 END
 END vss.gds78
 PIN vss.gds79
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 2.9235 12.818 3.1235 ;
 END
 END vss.gds79
 PIN vss.gds80
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 1.418 13.898 1.618 ;
 END
 END vss.gds80
 PIN vss.gds81
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 14 1.596 14.056 1.769 ;
 RECT 14.168 1.569 14.224 1.769 ;
 RECT 14.84 1.613 14.896 1.778 ;
 RECT 14 5.376 14.056 5.549 ;
 RECT 14.168 5.349 14.224 5.549 ;
 RECT 14 2.856 14.056 3.029 ;
 RECT 14.168 2.829 14.224 3.029 ;
 RECT 14 4.116 14.056 4.289 ;
 RECT 14.168 4.089 14.224 4.289 ;
 RECT 14.336 4.709 14.392 4.909 ;
 RECT 14.168 4.709 14.224 4.909 ;
 RECT 14.336 2.189 14.392 2.389 ;
 RECT 14.168 2.189 14.224 2.389 ;
 RECT 14.336 3.449 14.392 3.649 ;
 RECT 14.168 3.449 14.224 3.649 ;
 RECT 15.008 3.659 15.064 3.859 ;
 RECT 14.84 4.133 14.896 4.298 ;
 RECT 14.672 4.133 14.728 4.298 ;
 RECT 13.664 3.583 13.72 3.783 ;
 RECT 15.008 2.399 15.064 2.599 ;
 RECT 14.84 2.873 14.896 3.038 ;
 RECT 14.672 2.873 14.728 3.038 ;
 RECT 13.664 2.323 13.72 2.523 ;
 RECT 15.008 4.919 15.064 5.119 ;
 RECT 14.84 5.393 14.896 5.558 ;
 RECT 14.672 5.393 14.728 5.558 ;
 RECT 13.664 4.843 13.72 5.043 ;
 RECT 14.336 0.929 14.392 1.129 ;
 RECT 14.168 0.929 14.224 1.129 ;
 RECT 15.008 1.139 15.064 1.339 ;
 RECT 15.176 3.0995 15.232 3.2995 ;
 RECT 14.672 1.613 14.728 1.778 ;
 RECT 13.664 1.063 13.72 1.263 ;
 RECT 12.824 2.884 12.88 3.084 ;
 RECT 13.496 2.895 13.552 3.095 ;
 RECT 12.488 2.914 12.544 3.114 ;
 RECT 13.328 2.833 13.384 3.033 ;
 RECT 13.16 2.884 13.216 3.084 ;
 RECT 12.992 2.884 13.048 3.084 ;
 RECT 12.656 2.914 12.712 3.114 ;
 END
 END vss.gds81
 PIN vss.gds82
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 2.916 15.418 3.116 ;
 END
 END vss.gds82
 PIN vss.gds83
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 2.9095 20.274 3.1095 ;
 END
 END vss.gds83
 PIN vss.gds84
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 2.9095 18.93 3.1095 ;
 END
 END vss.gds84
 PIN vss.gds85
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.038 2.9095 19.098 3.1095 ;
 END
 END vss.gds85
 PIN vss.gds86
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.206 2.9095 19.266 3.1095 ;
 END
 END vss.gds86
 PIN vss.gds87
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.374 2.9095 19.434 3.1095 ;
 END
 END vss.gds87
 PIN vss.gds88
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 2.9095 19.602 3.1095 ;
 END
 END vss.gds88
 PIN vss.gds89
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 2.9235 17.314 3.1235 ;
 END
 END vss.gds89
 PIN vss.gds90
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 2.9785 16.994 3.1785 ;
 END
 END vss.gds90
 PIN vss.gds91
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.71 2.9095 19.77 3.1095 ;
 END
 END vss.gds91
 PIN vss.gds92
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.878 2.9095 19.938 3.1095 ;
 END
 END vss.gds92
 PIN vss.gds93
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 3.06 15.842 3.26 ;
 END
 END vss.gds93
 PIN vss.gds94
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 3.072 16.814 3.272 ;
 END
 END vss.gds94
 PIN vss.gds95
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 4.693 16.146 4.893 ;
 END
 END vss.gds95
 PIN vss.gds96
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.046 2.9095 20.106 3.1095 ;
 END
 END vss.gds96
 PIN vss.gds97
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.702 2.9095 18.762 3.1095 ;
 END
 END vss.gds97
 PIN vss.gds98
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.534 2.9095 18.594 3.1095 ;
 END
 END vss.gds98
 PIN vss.gds99
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.366 2.9095 18.426 3.1095 ;
 END
 END vss.gds99
 PIN vss.gds100
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 2.941 18.258 3.141 ;
 END
 END vss.gds100
 PIN vss.gds101
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 2.9235 17.834 3.1235 ;
 END
 END vss.gds101
 PIN vss.gds102
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 3.433 16.146 3.633 ;
 END
 END vss.gds102
 PIN vss.gds103
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 2.173 16.146 2.373 ;
 END
 END vss.gds103
 PIN vss.gds104
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 0.913 16.146 1.113 ;
 END
 END vss.gds104
 PIN vss.gds105
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.438 3.0755 17.494 3.2755 ;
 END
 END vss.gds105
 PIN vss.gds106
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 2.8265 16.49 3.0265 ;
 END
 END vss.gds106
 PIN vss.gds107
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.986 2.803 18.026 3.003 ;
 END
 END vss.gds107
 PIN vss.gds108
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 15.596 0.58 15.652 0.78 ;
 RECT 15.848 0.583 15.904 0.783 ;
 RECT 16.52 1.616 16.576 1.769 ;
 RECT 15.764 1.613 15.82 1.778 ;
 RECT 15.596 1.613 15.652 1.778 ;
 RECT 15.596 4.36 15.652 4.56 ;
 RECT 15.848 4.363 15.904 4.563 ;
 RECT 16.52 5.396 16.576 5.549 ;
 RECT 15.764 5.393 15.82 5.558 ;
 RECT 15.596 5.393 15.652 5.558 ;
 RECT 15.596 1.84 15.652 2.04 ;
 RECT 15.848 1.843 15.904 2.043 ;
 RECT 16.52 2.876 16.576 3.029 ;
 RECT 15.764 2.873 15.82 3.038 ;
 RECT 15.596 2.873 15.652 3.038 ;
 RECT 15.596 3.1 15.652 3.3 ;
 RECT 15.848 3.103 15.904 3.303 ;
 RECT 16.52 4.136 16.576 4.289 ;
 RECT 15.764 4.133 15.82 4.298 ;
 RECT 15.596 4.133 15.652 4.298 ;
 RECT 15.428 3.659 15.484 3.859 ;
 RECT 16.352 3.7595 16.408 3.9595 ;
 RECT 16.856 3.5075 16.912 3.7075 ;
 RECT 15.428 2.399 15.484 2.599 ;
 RECT 16.352 2.4995 16.408 2.6995 ;
 RECT 16.856 2.2475 16.912 2.4475 ;
 RECT 15.428 4.919 15.484 5.119 ;
 RECT 16.352 5.0195 16.408 5.2195 ;
 RECT 16.856 4.7675 16.912 4.9675 ;
 RECT 15.428 1.139 15.484 1.339 ;
 RECT 16.352 1.2395 16.408 1.4395 ;
 RECT 16.856 0.9875 16.912 1.1875 ;
 RECT 17.864 2.914 17.92 3.114 ;
 RECT 17.696 2.9215 17.752 3.1215 ;
 RECT 17.528 2.914 17.584 3.114 ;
 RECT 17.36 2.914 17.416 3.114 ;
 RECT 17.192 2.914 17.248 3.114 ;
 RECT 18.032 2.914 18.088 3.114 ;
 RECT 17.024 3.029 17.08 3.229 ;
 END
 END vss.gds108
 PIN vss.gds109
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.17 2.9095 25.23 3.1095 ;
 END
 END vss.gds109
 PIN vss.gds110
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.002 2.9095 25.062 3.1095 ;
 END
 END vss.gds110
 PIN vss.gds111
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.834 2.9095 24.894 3.1095 ;
 END
 END vss.gds111
 PIN vss.gds112
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.498 2.9095 24.558 3.1095 ;
 END
 END vss.gds112
 PIN vss.gds113
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.33 2.9095 24.39 3.1095 ;
 END
 END vss.gds113
 PIN vss.gds114
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.162 2.9095 24.222 3.1095 ;
 END
 END vss.gds114
 PIN vss.gds115
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.382 2.9095 20.442 3.1095 ;
 END
 END vss.gds115
 PIN vss.gds116
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.55 2.9095 20.61 3.1095 ;
 END
 END vss.gds116
 PIN vss.gds117
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.718 2.9095 20.778 3.1095 ;
 END
 END vss.gds117
 PIN vss.gds118
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.054 2.9095 21.114 3.1095 ;
 END
 END vss.gds118
 PIN vss.gds119
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.222 2.9095 21.282 3.1095 ;
 END
 END vss.gds119
 PIN vss.gds120
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.39 2.9095 21.45 3.1095 ;
 END
 END vss.gds120
 PIN vss.gds121
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.726 2.9095 21.786 3.1095 ;
 END
 END vss.gds121
 PIN vss.gds122
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.894 2.9095 21.954 3.1095 ;
 END
 END vss.gds122
 PIN vss.gds123
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.062 2.9095 22.122 3.1095 ;
 END
 END vss.gds123
 PIN vss.gds124
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.398 2.9095 22.458 3.1095 ;
 END
 END vss.gds124
 PIN vss.gds125
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.566 2.9095 22.626 3.1095 ;
 END
 END vss.gds125
 PIN vss.gds126
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.734 2.9095 22.794 3.1095 ;
 END
 END vss.gds126
 PIN vss.gds127
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 2.9095 24.726 3.1095 ;
 END
 END vss.gds127
 PIN vss.gds128
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 2.9095 21.618 3.1095 ;
 END
 END vss.gds128
 PIN vss.gds129
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 2.9095 20.946 3.1095 ;
 END
 END vss.gds129
 PIN vss.gds130
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 2.9095 22.29 3.1095 ;
 END
 END vss.gds130
 PIN vss.gds131
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 2.9095 22.962 3.1095 ;
 END
 END vss.gds131
 PIN vss.gds132
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.07 2.9095 23.13 3.1095 ;
 END
 END vss.gds132
 PIN vss.gds133
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.238 2.9095 23.298 3.1095 ;
 END
 END vss.gds133
 PIN vss.gds134
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.406 2.9095 23.466 3.1095 ;
 END
 END vss.gds134
 PIN vss.gds135
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 2.9095 23.634 3.1095 ;
 END
 END vss.gds135
 PIN vss.gds136
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 23.912 3.596 23.968 3.796 ;
 RECT 23.912 2.336 23.968 2.536 ;
 RECT 23.912 4.856 23.968 5.056 ;
 RECT 23.912 1.076 23.968 1.276 ;
 RECT 23.744 2.966 23.8 3.166 ;
 END
 END vss.gds136
 PIN vss.gds137
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.202 2.9095 29.262 3.1095 ;
 END
 END vss.gds137
 PIN vss.gds138
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.034 2.9095 29.094 3.1095 ;
 END
 END vss.gds138
 PIN vss.gds139
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.866 2.9095 28.926 3.1095 ;
 END
 END vss.gds139
 PIN vss.gds140
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.53 2.9095 28.59 3.1095 ;
 END
 END vss.gds140
 PIN vss.gds141
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.362 2.9095 28.422 3.1095 ;
 END
 END vss.gds141
 PIN vss.gds142
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.194 2.9095 28.254 3.1095 ;
 END
 END vss.gds142
 PIN vss.gds143
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.858 2.9095 27.918 3.1095 ;
 END
 END vss.gds143
 PIN vss.gds144
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.69 2.9095 27.75 3.1095 ;
 END
 END vss.gds144
 PIN vss.gds145
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.522 2.9095 27.582 3.1095 ;
 END
 END vss.gds145
 PIN vss.gds146
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.186 2.9095 27.246 3.1095 ;
 END
 END vss.gds146
 PIN vss.gds147
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.018 2.9095 27.078 3.1095 ;
 END
 END vss.gds147
 PIN vss.gds148
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.85 2.9095 26.91 3.1095 ;
 END
 END vss.gds148
 PIN vss.gds149
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.514 2.9095 26.574 3.1095 ;
 END
 END vss.gds149
 PIN vss.gds150
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.346 2.9095 26.406 3.1095 ;
 END
 END vss.gds150
 PIN vss.gds151
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.178 2.9095 26.238 3.1095 ;
 END
 END vss.gds151
 PIN vss.gds152
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.842 2.9095 25.902 3.1095 ;
 END
 END vss.gds152
 PIN vss.gds153
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.674 2.9095 25.734 3.1095 ;
 END
 END vss.gds153
 PIN vss.gds154
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.506 2.9095 25.566 3.1095 ;
 END
 END vss.gds154
 PIN vss.gds155
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 2.9095 28.758 3.1095 ;
 END
 END vss.gds155
 PIN vss.gds156
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 2.9095 28.086 3.1095 ;
 END
 END vss.gds156
 PIN vss.gds157
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 2.9095 27.414 3.1095 ;
 END
 END vss.gds157
 PIN vss.gds158
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 2.9095 26.742 3.1095 ;
 END
 END vss.gds158
 PIN vss.gds159
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 2.9095 26.07 3.1095 ;
 END
 END vss.gds159
 PIN vss.gds160
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 2.9095 25.398 3.1095 ;
 END
 END vss.gds160
 PIN vss.gds161
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 2.941 29.43 3.141 ;
 END
 END vss.gds161
 PIN vss.gds162
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 3.0755 30.11 3.2755 ;
 END
 END vss.gds162
 PIN vss.gds163
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 2.9235 29.87 3.1235 ;
 END
 END vss.gds163
 PIN vss.gds164
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 2.803 29.642 3.003 ;
 END
 END vss.gds164
 PIN vss.gds165
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.876 2.884 29.932 3.084 ;
 RECT 30.212 2.884 30.268 3.084 ;
 RECT 29.54 2.914 29.596 3.114 ;
 RECT 30.044 2.884 30.1 3.084 ;
 RECT 29.708 2.914 29.764 3.114 ;
 END
 END vss.gds165
 PIN vss.gds166
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 1.458 31.922 1.658 ;
 END
 END vss.gds166
 PIN vss.gds167
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 1.418 30.95 1.618 ;
 END
 END vss.gds167
 PIN vss.gds168
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 5.238 31.922 5.438 ;
 END
 END vss.gds168
 PIN vss.gds169
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 2.678 30.95 2.878 ;
 END
 END vss.gds169
 PIN vss.gds170
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 2.718 31.922 2.918 ;
 END
 END vss.gds170
 PIN vss.gds171
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 3.938 30.95 4.138 ;
 END
 END vss.gds171
 PIN vss.gds172
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 3.978 31.922 4.178 ;
 END
 END vss.gds172
 PIN vss.gds173
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.314 3.072 30.37 3.272 ;
 END
 END vss.gds173
 PIN vss.gds174
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 3.06 32.214 3.26 ;
 END
 END vss.gds174
 PIN vss.gds175
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 2.9785 34.046 3.1785 ;
 END
 END vss.gds175
 PIN vss.gds176
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 3.0195 30.71 3.2195 ;
 END
 END vss.gds176
 PIN vss.gds177
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 3.06 32.894 3.26 ;
 END
 END vss.gds177
 PIN vss.gds178
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 2.8265 33.542 3.0265 ;
 END
 END vss.gds178
 PIN vss.gds179
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 3.06 31.55 3.26 ;
 END
 END vss.gds179
 PIN vss.gds180
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 3.072 33.866 3.272 ;
 END
 END vss.gds180
 PIN vss.gds181
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 2.9235 34.886 3.1235 ;
 END
 END vss.gds181
 PIN vss.gds182
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.49 3.0755 34.546 3.2755 ;
 END
 END vss.gds182
 PIN vss.gds183
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 2.916 32.47 3.116 ;
 END
 END vss.gds183
 PIN vss.gds184
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 4.693 33.198 4.893 ;
 END
 END vss.gds184
 PIN vss.gds185
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 3.433 33.198 3.633 ;
 END
 END vss.gds185
 PIN vss.gds186
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 2.173 33.198 2.373 ;
 END
 END vss.gds186
 PIN vss.gds187
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 0.913 33.198 1.113 ;
 END
 END vss.gds187
 PIN vss.gds188
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 5.198 30.95 5.398 ;
 END
 END vss.gds188
 PIN vss.gds189
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 2.9235 34.366 3.1235 ;
 END
 END vss.gds189
 PIN vss.gds190
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.038 2.803 35.078 3.003 ;
 END
 END vss.gds190
 PIN vss.gds191
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 32.648 0.58 32.704 0.78 ;
 RECT 32.9 0.583 32.956 0.783 ;
 RECT 33.572 1.616 33.628 1.769 ;
 RECT 31.052 1.596 31.108 1.769 ;
 RECT 31.22 1.569 31.276 1.769 ;
 RECT 32.816 1.613 32.872 1.778 ;
 RECT 32.648 1.613 32.704 1.778 ;
 RECT 31.892 1.613 31.948 1.778 ;
 RECT 31.724 1.613 31.78 1.778 ;
 RECT 31.388 0.929 31.444 1.129 ;
 RECT 31.22 0.929 31.276 1.129 ;
 RECT 30.716 1.063 30.772 1.263 ;
 RECT 32.648 4.36 32.704 4.56 ;
 RECT 32.9 4.363 32.956 4.563 ;
 RECT 33.572 5.396 33.628 5.549 ;
 RECT 31.052 5.376 31.108 5.549 ;
 RECT 31.22 5.349 31.276 5.549 ;
 RECT 32.816 5.393 32.872 5.558 ;
 RECT 32.648 5.393 32.704 5.558 ;
 RECT 31.892 5.393 31.948 5.558 ;
 RECT 31.724 5.393 31.78 5.558 ;
 RECT 32.648 1.84 32.704 2.04 ;
 RECT 32.9 1.843 32.956 2.043 ;
 RECT 33.572 2.876 33.628 3.029 ;
 RECT 31.052 2.856 31.108 3.029 ;
 RECT 31.22 2.829 31.276 3.029 ;
 RECT 32.816 2.873 32.872 3.038 ;
 RECT 32.648 2.873 32.704 3.038 ;
 RECT 31.892 2.873 31.948 3.038 ;
 RECT 31.724 2.873 31.78 3.038 ;
 RECT 33.572 4.136 33.628 4.289 ;
 RECT 31.052 4.116 31.108 4.289 ;
 RECT 31.22 4.089 31.276 4.289 ;
 RECT 32.816 4.133 32.872 4.298 ;
 RECT 32.648 4.133 32.704 4.298 ;
 RECT 31.892 4.133 31.948 4.298 ;
 RECT 31.724 4.133 31.78 4.298 ;
 RECT 32.648 3.1 32.704 3.3 ;
 RECT 32.9 3.103 32.956 3.303 ;
 RECT 31.388 2.189 31.444 2.389 ;
 RECT 31.22 2.189 31.276 2.389 ;
 RECT 31.388 4.709 31.444 4.909 ;
 RECT 31.22 4.709 31.276 4.909 ;
 RECT 32.06 4.919 32.116 5.119 ;
 RECT 32.48 4.919 32.536 5.119 ;
 RECT 32.06 1.139 32.116 1.339 ;
 RECT 32.48 1.139 32.536 1.339 ;
 RECT 31.388 3.449 31.444 3.649 ;
 RECT 31.22 3.449 31.276 3.649 ;
 RECT 33.404 3.7595 33.46 3.9595 ;
 RECT 33.908 3.5075 33.964 3.7075 ;
 RECT 30.716 2.323 30.772 2.523 ;
 RECT 32.06 2.399 32.116 2.599 ;
 RECT 32.48 2.399 32.536 2.599 ;
 RECT 30.716 3.583 30.772 3.783 ;
 RECT 32.06 3.659 32.116 3.859 ;
 RECT 32.48 3.659 32.536 3.859 ;
 RECT 30.716 4.843 30.772 5.043 ;
 RECT 33.404 5.0195 33.46 5.2195 ;
 RECT 33.908 4.7675 33.964 4.9675 ;
 RECT 30.548 2.895 30.604 3.095 ;
 RECT 33.404 2.4995 33.46 2.6995 ;
 RECT 33.908 2.2475 33.964 2.4475 ;
 RECT 30.38 2.833 30.436 3.033 ;
 RECT 32.228 3.0995 32.284 3.2995 ;
 RECT 33.404 1.2395 33.46 1.4395 ;
 RECT 33.908 0.9875 33.964 1.1875 ;
 RECT 34.916 2.914 34.972 3.114 ;
 RECT 34.748 2.9215 34.804 3.1215 ;
 RECT 34.58 2.914 34.636 3.114 ;
 RECT 34.412 2.914 34.468 3.114 ;
 RECT 34.244 2.914 34.3 3.114 ;
 RECT 35.084 2.914 35.14 3.114 ;
 RECT 34.076 3.029 34.132 3.229 ;
 END
 END vss.gds191
 PIN vss.gds192
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.122 2.9095 40.182 3.1095 ;
 END
 END vss.gds192
 PIN vss.gds193
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.754 2.9095 35.814 3.1095 ;
 END
 END vss.gds193
 PIN vss.gds194
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.09 2.9095 36.15 3.1095 ;
 END
 END vss.gds194
 PIN vss.gds195
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.258 2.9095 36.318 3.1095 ;
 END
 END vss.gds195
 PIN vss.gds196
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.426 2.9095 36.486 3.1095 ;
 END
 END vss.gds196
 PIN vss.gds197
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.762 2.9095 36.822 3.1095 ;
 END
 END vss.gds197
 PIN vss.gds198
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.93 2.9095 36.99 3.1095 ;
 END
 END vss.gds198
 PIN vss.gds199
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.098 2.9095 37.158 3.1095 ;
 END
 END vss.gds199
 PIN vss.gds200
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.434 2.9095 37.494 3.1095 ;
 END
 END vss.gds200
 PIN vss.gds201
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.602 2.9095 37.662 3.1095 ;
 END
 END vss.gds201
 PIN vss.gds202
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.77 2.9095 37.83 3.1095 ;
 END
 END vss.gds202
 PIN vss.gds203
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.106 2.9095 38.166 3.1095 ;
 END
 END vss.gds203
 PIN vss.gds204
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.274 2.9095 38.334 3.1095 ;
 END
 END vss.gds204
 PIN vss.gds205
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 2.9095 36.654 3.1095 ;
 END
 END vss.gds205
 PIN vss.gds206
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 2.9095 37.326 3.1095 ;
 END
 END vss.gds206
 PIN vss.gds207
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 2.9095 37.998 3.1095 ;
 END
 END vss.gds207
 PIN vss.gds208
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.442 2.9095 38.502 3.1095 ;
 END
 END vss.gds208
 PIN vss.gds209
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 2.9095 38.67 3.1095 ;
 END
 END vss.gds209
 PIN vss.gds210
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.778 2.9095 38.838 3.1095 ;
 END
 END vss.gds210
 PIN vss.gds211
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 2.9095 35.982 3.1095 ;
 END
 END vss.gds211
 PIN vss.gds212
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.946 2.9095 39.006 3.1095 ;
 END
 END vss.gds212
 PIN vss.gds213
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.586 2.9095 35.646 3.1095 ;
 END
 END vss.gds213
 PIN vss.gds214
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.45 2.9095 39.51 3.1095 ;
 END
 END vss.gds214
 PIN vss.gds215
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.618 2.9095 39.678 3.1095 ;
 END
 END vss.gds215
 PIN vss.gds216
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.114 2.9095 39.174 3.1095 ;
 END
 END vss.gds216
 PIN vss.gds217
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.786 2.9095 39.846 3.1095 ;
 END
 END vss.gds217
 PIN vss.gds218
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 2.9095 40.014 3.1095 ;
 END
 END vss.gds218
 PIN vss.gds219
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.418 2.9095 35.478 3.1095 ;
 END
 END vss.gds219
 PIN vss.gds220
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 2.941 35.31 3.141 ;
 END
 END vss.gds220
 PIN vss.gds221
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 2.9095 39.342 3.1095 ;
 END
 END vss.gds221
 PIN vss.gds222
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.91 2.9095 44.97 3.1095 ;
 END
 END vss.gds222
 PIN vss.gds223
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.742 2.9095 44.802 3.1095 ;
 END
 END vss.gds223
 PIN vss.gds224
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.574 2.9095 44.634 3.1095 ;
 END
 END vss.gds224
 PIN vss.gds225
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.238 2.9095 44.298 3.1095 ;
 END
 END vss.gds225
 PIN vss.gds226
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.07 2.9095 44.13 3.1095 ;
 END
 END vss.gds226
 PIN vss.gds227
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.902 2.9095 43.962 3.1095 ;
 END
 END vss.gds227
 PIN vss.gds228
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.566 2.9095 43.626 3.1095 ;
 END
 END vss.gds228
 PIN vss.gds229
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.398 2.9095 43.458 3.1095 ;
 END
 END vss.gds229
 PIN vss.gds230
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.23 2.9095 43.29 3.1095 ;
 END
 END vss.gds230
 PIN vss.gds231
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.894 2.9095 42.954 3.1095 ;
 END
 END vss.gds231
 PIN vss.gds232
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.726 2.9095 42.786 3.1095 ;
 END
 END vss.gds232
 PIN vss.gds233
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.558 2.9095 42.618 3.1095 ;
 END
 END vss.gds233
 PIN vss.gds234
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.222 2.9095 42.282 3.1095 ;
 END
 END vss.gds234
 PIN vss.gds235
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.054 2.9095 42.114 3.1095 ;
 END
 END vss.gds235
 PIN vss.gds236
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.886 2.9095 41.946 3.1095 ;
 END
 END vss.gds236
 PIN vss.gds237
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.55 2.9095 41.61 3.1095 ;
 END
 END vss.gds237
 PIN vss.gds238
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.382 2.9095 41.442 3.1095 ;
 END
 END vss.gds238
 PIN vss.gds239
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.214 2.9095 41.274 3.1095 ;
 END
 END vss.gds239
 PIN vss.gds240
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.29 2.9095 40.35 3.1095 ;
 END
 END vss.gds240
 PIN vss.gds241
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.458 2.9095 40.518 3.1095 ;
 END
 END vss.gds241
 PIN vss.gds242
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 2.9095 45.138 3.1095 ;
 END
 END vss.gds242
 PIN vss.gds243
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 2.9095 44.466 3.1095 ;
 END
 END vss.gds243
 PIN vss.gds244
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 2.9095 43.794 3.1095 ;
 END
 END vss.gds244
 PIN vss.gds245
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 2.9095 43.122 3.1095 ;
 END
 END vss.gds245
 PIN vss.gds246
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 2.9095 42.45 3.1095 ;
 END
 END vss.gds246
 PIN vss.gds247
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 2.9095 41.778 3.1095 ;
 END
 END vss.gds247
 PIN vss.gds248
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 2.9095 40.686 3.1095 ;
 END
 END vss.gds248
 PIN vss.gds249
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 40.964 4.856 41.02 5.056 ;
 RECT 40.964 3.596 41.02 3.796 ;
 RECT 40.964 2.336 41.02 2.536 ;
 RECT 40.964 1.076 41.02 1.276 ;
 RECT 40.796 2.966 40.852 3.166 ;
 END
 END vss.gds249
 PIN vss.gds250
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 1.458 48.974 1.658 ;
 END
 END vss.gds250
 PIN vss.gds251
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 1.418 48.002 1.618 ;
 END
 END vss.gds251
 PIN vss.gds252
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 5.238 48.974 5.438 ;
 END
 END vss.gds252
 PIN vss.gds253
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 2.718 48.974 2.918 ;
 END
 END vss.gds253
 PIN vss.gds254
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 3.978 48.974 4.178 ;
 END
 END vss.gds254
 PIN vss.gds255
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 3.938 48.002 4.138 ;
 END
 END vss.gds255
 PIN vss.gds256
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 5.198 48.002 5.398 ;
 END
 END vss.gds256
 PIN vss.gds257
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.366 3.072 47.422 3.272 ;
 END
 END vss.gds257
 PIN vss.gds258
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.254 2.9095 46.314 3.1095 ;
 END
 END vss.gds258
 PIN vss.gds259
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.086 2.9095 46.146 3.1095 ;
 END
 END vss.gds259
 PIN vss.gds260
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.918 2.9095 45.978 3.1095 ;
 END
 END vss.gds260
 PIN vss.gds261
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.582 2.9095 45.642 3.1095 ;
 END
 END vss.gds261
 PIN vss.gds262
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.414 2.9095 45.474 3.1095 ;
 END
 END vss.gds262
 PIN vss.gds263
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.246 2.9095 45.306 3.1095 ;
 END
 END vss.gds263
 PIN vss.gds264
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 3.0755 47.162 3.2755 ;
 END
 END vss.gds264
 PIN vss.gds265
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 2.941 46.482 3.141 ;
 END
 END vss.gds265
 PIN vss.gds266
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 2.9095 45.81 3.1095 ;
 END
 END vss.gds266
 PIN vss.gds267
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 2.9235 46.922 3.1235 ;
 END
 END vss.gds267
 PIN vss.gds268
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 2.803 46.694 3.003 ;
 END
 END vss.gds268
 PIN vss.gds269
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 3.0195 47.762 3.2195 ;
 END
 END vss.gds269
 PIN vss.gds270
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 3.06 49.266 3.26 ;
 END
 END vss.gds270
 PIN vss.gds271
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 3.06 48.602 3.26 ;
 END
 END vss.gds271
 PIN vss.gds272
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 3.06 49.946 3.26 ;
 END
 END vss.gds272
 PIN vss.gds273
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 4.693 50.25 4.893 ;
 END
 END vss.gds273
 PIN vss.gds274
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 3.433 50.25 3.633 ;
 END
 END vss.gds274
 PIN vss.gds275
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 2.173 50.25 2.373 ;
 END
 END vss.gds275
 PIN vss.gds276
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 0.913 50.25 1.113 ;
 END
 END vss.gds276
 PIN vss.gds277
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 2.916 49.522 3.116 ;
 END
 END vss.gds277
 PIN vss.gds278
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 2.678 48.002 2.878 ;
 END
 END vss.gds278
 PIN vss.gds279
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 48.104 1.596 48.16 1.769 ;
 RECT 48.272 1.569 48.328 1.769 ;
 RECT 49.868 1.613 49.924 1.778 ;
 RECT 49.7 1.613 49.756 1.778 ;
 RECT 48.944 1.613 49 1.778 ;
 RECT 48.776 1.613 48.832 1.778 ;
 RECT 49.7 0.58 49.756 0.78 ;
 RECT 49.952 0.583 50.008 0.783 ;
 RECT 48.44 0.929 48.496 1.129 ;
 RECT 48.272 0.929 48.328 1.129 ;
 RECT 47.768 1.063 47.824 1.263 ;
 RECT 49.7 1.84 49.756 2.04 ;
 RECT 49.952 1.843 50.008 2.043 ;
 RECT 49.7 4.36 49.756 4.56 ;
 RECT 49.952 4.363 50.008 4.563 ;
 RECT 48.104 5.376 48.16 5.549 ;
 RECT 48.272 5.349 48.328 5.549 ;
 RECT 49.868 5.393 49.924 5.558 ;
 RECT 49.7 5.393 49.756 5.558 ;
 RECT 48.944 5.393 49 5.558 ;
 RECT 48.776 5.393 48.832 5.558 ;
 RECT 48.104 2.856 48.16 3.029 ;
 RECT 48.272 2.829 48.328 3.029 ;
 RECT 49.868 2.873 49.924 3.038 ;
 RECT 49.7 2.873 49.756 3.038 ;
 RECT 48.944 2.873 49 3.038 ;
 RECT 48.776 2.873 48.832 3.038 ;
 RECT 48.104 4.116 48.16 4.289 ;
 RECT 48.272 4.089 48.328 4.289 ;
 RECT 49.868 4.133 49.924 4.298 ;
 RECT 49.7 4.133 49.756 4.298 ;
 RECT 48.944 4.133 49 4.298 ;
 RECT 48.776 4.133 48.832 4.298 ;
 RECT 49.7 3.1 49.756 3.3 ;
 RECT 49.952 3.103 50.008 3.303 ;
 RECT 48.44 4.709 48.496 4.909 ;
 RECT 48.272 4.709 48.328 4.909 ;
 RECT 47.768 4.843 47.824 5.043 ;
 RECT 49.112 4.919 49.168 5.119 ;
 RECT 49.532 4.919 49.588 5.119 ;
 RECT 48.44 3.449 48.496 3.649 ;
 RECT 48.272 3.449 48.328 3.649 ;
 RECT 47.768 3.583 47.824 3.783 ;
 RECT 49.112 3.659 49.168 3.859 ;
 RECT 49.532 3.659 49.588 3.859 ;
 RECT 49.112 1.139 49.168 1.339 ;
 RECT 49.532 1.139 49.588 1.339 ;
 RECT 48.44 2.189 48.496 2.389 ;
 RECT 48.272 2.189 48.328 2.389 ;
 RECT 49.112 2.399 49.168 2.599 ;
 RECT 49.532 2.399 49.588 2.599 ;
 RECT 47.768 2.323 47.824 2.523 ;
 RECT 47.6 2.895 47.656 3.095 ;
 RECT 47.432 2.833 47.488 3.033 ;
 RECT 47.264 2.884 47.32 3.084 ;
 RECT 46.928 2.884 46.984 3.084 ;
 RECT 47.096 2.884 47.152 3.084 ;
 RECT 49.28 3.0995 49.336 3.2995 ;
 RECT 46.592 2.914 46.648 3.114 ;
 RECT 46.76 2.914 46.816 3.114 ;
 END
 END vss.gds279
 PIN vss.gds280
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.638 2.9095 52.698 3.1095 ;
 END
 END vss.gds280
 PIN vss.gds281
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.806 2.9095 52.866 3.1095 ;
 END
 END vss.gds281
 PIN vss.gds282
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.142 2.9095 53.202 3.1095 ;
 END
 END vss.gds282
 PIN vss.gds283
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.31 2.9095 53.37 3.1095 ;
 END
 END vss.gds283
 PIN vss.gds284
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.478 2.9095 53.538 3.1095 ;
 END
 END vss.gds284
 PIN vss.gds285
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.814 2.9095 53.874 3.1095 ;
 END
 END vss.gds285
 PIN vss.gds286
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.982 2.9095 54.042 3.1095 ;
 END
 END vss.gds286
 PIN vss.gds287
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.15 2.9095 54.21 3.1095 ;
 END
 END vss.gds287
 PIN vss.gds288
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.486 2.9095 54.546 3.1095 ;
 END
 END vss.gds288
 PIN vss.gds289
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.654 2.9095 54.714 3.1095 ;
 END
 END vss.gds289
 PIN vss.gds290
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.822 2.9095 54.882 3.1095 ;
 END
 END vss.gds290
 PIN vss.gds291
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.158 2.9095 55.218 3.1095 ;
 END
 END vss.gds291
 PIN vss.gds292
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 2.9095 55.05 3.1095 ;
 END
 END vss.gds292
 PIN vss.gds293
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 2.9095 54.378 3.1095 ;
 END
 END vss.gds293
 PIN vss.gds294
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 3.072 50.918 3.272 ;
 END
 END vss.gds294
 PIN vss.gds295
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 2.9095 53.706 3.1095 ;
 END
 END vss.gds295
 PIN vss.gds296
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 2.9785 51.098 3.1785 ;
 END
 END vss.gds296
 PIN vss.gds297
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 2.9095 53.034 3.1095 ;
 END
 END vss.gds297
 PIN vss.gds298
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 2.9235 51.938 3.1235 ;
 END
 END vss.gds298
 PIN vss.gds299
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.542 3.0755 51.598 3.2755 ;
 END
 END vss.gds299
 PIN vss.gds300
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 2.9235 51.418 3.1235 ;
 END
 END vss.gds300
 PIN vss.gds301
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 2.8265 50.594 3.0265 ;
 END
 END vss.gds301
 PIN vss.gds302
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.09 2.803 52.13 3.003 ;
 END
 END vss.gds302
 PIN vss.gds303
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.47 2.9095 52.53 3.1095 ;
 END
 END vss.gds303
 PIN vss.gds304
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 2.941 52.362 3.141 ;
 END
 END vss.gds304
 PIN vss.gds305
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 50.624 1.616 50.68 1.769 ;
 RECT 50.624 5.396 50.68 5.549 ;
 RECT 50.624 2.876 50.68 3.029 ;
 RECT 50.624 4.136 50.68 4.289 ;
 RECT 50.456 5.0195 50.512 5.2195 ;
 RECT 50.96 4.7675 51.016 4.9675 ;
 RECT 50.456 3.7595 50.512 3.9595 ;
 RECT 50.96 3.5075 51.016 3.7075 ;
 RECT 50.456 2.4995 50.512 2.6995 ;
 RECT 50.96 2.2475 51.016 2.4475 ;
 RECT 50.456 1.2395 50.512 1.4395 ;
 RECT 50.96 0.9875 51.016 1.1875 ;
 RECT 51.968 2.914 52.024 3.114 ;
 RECT 51.8 2.9215 51.856 3.1215 ;
 RECT 51.632 2.914 51.688 3.114 ;
 RECT 51.464 2.914 51.52 3.114 ;
 RECT 51.296 2.914 51.352 3.114 ;
 RECT 52.136 2.914 52.192 3.114 ;
 RECT 51.128 3.029 51.184 3.229 ;
 END
 END vss.gds305
 PIN vss.gds306
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.946 2.9095 60.006 3.1095 ;
 END
 END vss.gds306
 PIN vss.gds307
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.778 2.9095 59.838 3.1095 ;
 END
 END vss.gds307
 PIN vss.gds308
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.61 2.9095 59.67 3.1095 ;
 END
 END vss.gds308
 PIN vss.gds309
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.274 2.9095 59.334 3.1095 ;
 END
 END vss.gds309
 PIN vss.gds310
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.106 2.9095 59.166 3.1095 ;
 END
 END vss.gds310
 PIN vss.gds311
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.938 2.9095 58.998 3.1095 ;
 END
 END vss.gds311
 PIN vss.gds312
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.602 2.9095 58.662 3.1095 ;
 END
 END vss.gds312
 PIN vss.gds313
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.434 2.9095 58.494 3.1095 ;
 END
 END vss.gds313
 PIN vss.gds314
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.266 2.9095 58.326 3.1095 ;
 END
 END vss.gds314
 PIN vss.gds315
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.326 2.9095 55.386 3.1095 ;
 END
 END vss.gds315
 PIN vss.gds316
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.494 2.9095 55.554 3.1095 ;
 END
 END vss.gds316
 PIN vss.gds317
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 2.9095 60.174 3.1095 ;
 END
 END vss.gds317
 PIN vss.gds318
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 2.9095 59.502 3.1095 ;
 END
 END vss.gds318
 PIN vss.gds319
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 2.9095 58.83 3.1095 ;
 END
 END vss.gds319
 PIN vss.gds320
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 2.9095 55.722 3.1095 ;
 END
 END vss.gds320
 PIN vss.gds321
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.83 2.9095 55.89 3.1095 ;
 END
 END vss.gds321
 PIN vss.gds322
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.998 2.9095 56.058 3.1095 ;
 END
 END vss.gds322
 PIN vss.gds323
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.166 2.9095 56.226 3.1095 ;
 END
 END vss.gds323
 PIN vss.gds324
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 2.9095 56.394 3.1095 ;
 END
 END vss.gds324
 PIN vss.gds325
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.502 2.9095 56.562 3.1095 ;
 END
 END vss.gds325
 PIN vss.gds326
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.67 2.9095 56.73 3.1095 ;
 END
 END vss.gds326
 PIN vss.gds327
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.838 2.9095 56.898 3.1095 ;
 END
 END vss.gds327
 PIN vss.gds328
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.342 2.9095 57.402 3.1095 ;
 END
 END vss.gds328
 PIN vss.gds329
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.51 2.9095 57.57 3.1095 ;
 END
 END vss.gds329
 PIN vss.gds330
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 2.9095 57.738 3.1095 ;
 END
 END vss.gds330
 PIN vss.gds331
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.174 2.9095 57.234 3.1095 ;
 END
 END vss.gds331
 PIN vss.gds332
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 2.9095 57.066 3.1095 ;
 END
 END vss.gds332
 PIN vss.gds333
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 58.016 4.856 58.072 5.056 ;
 RECT 58.016 3.596 58.072 3.796 ;
 RECT 58.016 2.336 58.072 2.536 ;
 RECT 58.016 1.076 58.072 1.276 ;
 RECT 57.848 2.966 57.904 3.166 ;
 END
 END vss.gds333
 PIN vss.gds334
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 1.418 65.054 1.618 ;
 END
 END vss.gds334
 PIN vss.gds335
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 3.938 65.054 4.138 ;
 END
 END vss.gds335
 PIN vss.gds336
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 5.198 65.054 5.398 ;
 END
 END vss.gds336
 PIN vss.gds337
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 3.0755 64.214 3.2755 ;
 END
 END vss.gds337
 PIN vss.gds338
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.418 3.072 64.474 3.272 ;
 END
 END vss.gds338
 PIN vss.gds339
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.306 2.9095 63.366 3.1095 ;
 END
 END vss.gds339
 PIN vss.gds340
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.138 2.9095 63.198 3.1095 ;
 END
 END vss.gds340
 PIN vss.gds341
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.97 2.9095 63.03 3.1095 ;
 END
 END vss.gds341
 PIN vss.gds342
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.634 2.9095 62.694 3.1095 ;
 END
 END vss.gds342
 PIN vss.gds343
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.466 2.9095 62.526 3.1095 ;
 END
 END vss.gds343
 PIN vss.gds344
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.298 2.9095 62.358 3.1095 ;
 END
 END vss.gds344
 PIN vss.gds345
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.962 2.9095 62.022 3.1095 ;
 END
 END vss.gds345
 PIN vss.gds346
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.794 2.9095 61.854 3.1095 ;
 END
 END vss.gds346
 PIN vss.gds347
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.626 2.9095 61.686 3.1095 ;
 END
 END vss.gds347
 PIN vss.gds348
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.29 2.9095 61.35 3.1095 ;
 END
 END vss.gds348
 PIN vss.gds349
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.122 2.9095 61.182 3.1095 ;
 END
 END vss.gds349
 PIN vss.gds350
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.954 2.9095 61.014 3.1095 ;
 END
 END vss.gds350
 PIN vss.gds351
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.618 2.9095 60.678 3.1095 ;
 END
 END vss.gds351
 PIN vss.gds352
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.45 2.9095 60.51 3.1095 ;
 END
 END vss.gds352
 PIN vss.gds353
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.282 2.9095 60.342 3.1095 ;
 END
 END vss.gds353
 PIN vss.gds354
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 2.941 63.534 3.141 ;
 END
 END vss.gds354
 PIN vss.gds355
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 2.9095 62.862 3.1095 ;
 END
 END vss.gds355
 PIN vss.gds356
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 2.9095 62.19 3.1095 ;
 END
 END vss.gds356
 PIN vss.gds357
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 2.9095 61.518 3.1095 ;
 END
 END vss.gds357
 PIN vss.gds358
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 2.9095 60.846 3.1095 ;
 END
 END vss.gds358
 PIN vss.gds359
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 2.9235 63.974 3.1235 ;
 END
 END vss.gds359
 PIN vss.gds360
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 2.803 63.746 3.003 ;
 END
 END vss.gds360
 PIN vss.gds361
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 3.0195 64.814 3.2195 ;
 END
 END vss.gds361
 PIN vss.gds362
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 2.678 65.054 2.878 ;
 END
 END vss.gds362
 PIN vss.gds363
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 65.156 1.596 65.212 1.769 ;
 RECT 65.156 5.376 65.212 5.549 ;
 RECT 65.156 2.856 65.212 3.029 ;
 RECT 65.156 4.116 65.212 4.289 ;
 RECT 64.82 1.063 64.876 1.263 ;
 RECT 64.82 4.843 64.876 5.043 ;
 RECT 64.82 3.583 64.876 3.783 ;
 RECT 64.82 2.323 64.876 2.523 ;
 RECT 64.652 2.895 64.708 3.095 ;
 RECT 64.484 2.833 64.54 3.033 ;
 RECT 64.316 2.884 64.372 3.084 ;
 RECT 64.148 2.884 64.204 3.084 ;
 RECT 63.98 2.884 64.036 3.084 ;
 RECT 63.644 2.914 63.7 3.114 ;
 RECT 63.812 2.914 63.868 3.114 ;
 END
 END vss.gds363
 PIN vss.gds364
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 1.458 66.026 1.658 ;
 END
 END vss.gds364
 PIN vss.gds365
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 5.238 66.026 5.438 ;
 END
 END vss.gds365
 PIN vss.gds366
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 2.718 66.026 2.918 ;
 END
 END vss.gds366
 PIN vss.gds367
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 3.978 66.026 4.178 ;
 END
 END vss.gds367
 PIN vss.gds368
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 4.693 67.302 4.893 ;
 END
 END vss.gds368
 PIN vss.gds369
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.69 2.9095 69.75 3.1095 ;
 END
 END vss.gds369
 PIN vss.gds370
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.858 2.9095 69.918 3.1095 ;
 END
 END vss.gds370
 PIN vss.gds371
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.194 2.9095 70.254 3.1095 ;
 END
 END vss.gds371
 PIN vss.gds372
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 2.9785 68.15 3.1785 ;
 END
 END vss.gds372
 PIN vss.gds373
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 3.06 66.318 3.26 ;
 END
 END vss.gds373
 PIN vss.gds374
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 2.9095 70.086 3.1095 ;
 END
 END vss.gds374
 PIN vss.gds375
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 3.06 66.998 3.26 ;
 END
 END vss.gds375
 PIN vss.gds376
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 3.06 65.654 3.26 ;
 END
 END vss.gds376
 PIN vss.gds377
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 2.8265 67.646 3.0265 ;
 END
 END vss.gds377
 PIN vss.gds378
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 2.916 66.574 3.116 ;
 END
 END vss.gds378
 PIN vss.gds379
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 3.072 67.97 3.272 ;
 END
 END vss.gds379
 PIN vss.gds380
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 2.9235 68.99 3.1235 ;
 END
 END vss.gds380
 PIN vss.gds381
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 3.433 67.302 3.633 ;
 END
 END vss.gds381
 PIN vss.gds382
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 2.173 67.302 2.373 ;
 END
 END vss.gds382
 PIN vss.gds383
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 0.913 67.302 1.113 ;
 END
 END vss.gds383
 PIN vss.gds384
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.594 3.0755 68.65 3.2755 ;
 END
 END vss.gds384
 PIN vss.gds385
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 2.9235 68.47 3.1235 ;
 END
 END vss.gds385
 PIN vss.gds386
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.142 2.803 69.182 3.003 ;
 END
 END vss.gds386
 PIN vss.gds387
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.522 2.9095 69.582 3.1095 ;
 END
 END vss.gds387
 PIN vss.gds388
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 2.941 69.414 3.141 ;
 END
 END vss.gds388
 PIN vss.gds389
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 67.676 1.616 67.732 1.769 ;
 RECT 65.324 1.569 65.38 1.769 ;
 RECT 66.92 1.613 66.976 1.778 ;
 RECT 66.752 1.613 66.808 1.778 ;
 RECT 65.996 1.613 66.052 1.778 ;
 RECT 65.828 1.613 65.884 1.778 ;
 RECT 66.752 0.58 66.808 0.78 ;
 RECT 67.004 0.583 67.06 0.783 ;
 RECT 67.676 5.396 67.732 5.549 ;
 RECT 65.324 5.349 65.38 5.549 ;
 RECT 66.92 5.393 66.976 5.558 ;
 RECT 66.752 5.393 66.808 5.558 ;
 RECT 65.996 5.393 66.052 5.558 ;
 RECT 65.828 5.393 65.884 5.558 ;
 RECT 67.676 2.876 67.732 3.029 ;
 RECT 65.324 2.829 65.38 3.029 ;
 RECT 66.92 2.873 66.976 3.038 ;
 RECT 66.752 2.873 66.808 3.038 ;
 RECT 65.996 2.873 66.052 3.038 ;
 RECT 65.828 2.873 65.884 3.038 ;
 RECT 67.676 4.136 67.732 4.289 ;
 RECT 65.324 4.089 65.38 4.289 ;
 RECT 66.92 4.133 66.976 4.298 ;
 RECT 66.752 4.133 66.808 4.298 ;
 RECT 65.996 4.133 66.052 4.298 ;
 RECT 65.828 4.133 65.884 4.298 ;
 RECT 66.752 1.84 66.808 2.04 ;
 RECT 67.004 1.843 67.06 2.043 ;
 RECT 65.492 0.929 65.548 1.129 ;
 RECT 65.324 0.929 65.38 1.129 ;
 RECT 66.752 3.1 66.808 3.3 ;
 RECT 67.004 3.103 67.06 3.303 ;
 RECT 66.752 4.36 66.808 4.56 ;
 RECT 67.004 4.363 67.06 4.563 ;
 RECT 65.492 4.709 65.548 4.909 ;
 RECT 65.324 4.709 65.38 4.909 ;
 RECT 68.012 4.7675 68.068 4.9675 ;
 RECT 67.508 5.0195 67.564 5.2195 ;
 RECT 67.508 3.7595 67.564 3.9595 ;
 RECT 68.012 3.5075 68.068 3.7075 ;
 RECT 65.492 3.449 65.548 3.649 ;
 RECT 65.324 3.449 65.38 3.649 ;
 RECT 66.164 1.139 66.22 1.339 ;
 RECT 66.584 1.139 66.64 1.339 ;
 RECT 65.492 2.189 65.548 2.389 ;
 RECT 65.324 2.189 65.38 2.389 ;
 RECT 66.164 2.399 66.22 2.599 ;
 RECT 66.584 2.399 66.64 2.599 ;
 RECT 66.164 4.919 66.22 5.119 ;
 RECT 66.584 4.919 66.64 5.119 ;
 RECT 66.164 3.659 66.22 3.859 ;
 RECT 66.584 3.659 66.64 3.859 ;
 RECT 67.508 2.4995 67.564 2.6995 ;
 RECT 68.012 2.2475 68.068 2.4475 ;
 RECT 68.012 0.9875 68.068 1.1875 ;
 RECT 67.508 1.2395 67.564 1.4395 ;
 RECT 66.332 3.0995 66.388 3.2995 ;
 RECT 69.02 2.914 69.076 3.114 ;
 RECT 68.852 2.9215 68.908 3.1215 ;
 RECT 68.684 2.914 68.74 3.114 ;
 RECT 68.516 2.914 68.572 3.114 ;
 RECT 68.348 2.914 68.404 3.114 ;
 RECT 69.188 2.914 69.244 3.114 ;
 RECT 68.18 3.029 68.236 3.229 ;
 END
 END vss.gds389
 PIN vss.gds390
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.362 2.9095 70.422 3.1095 ;
 END
 END vss.gds390
 PIN vss.gds391
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.53 2.9095 70.59 3.1095 ;
 END
 END vss.gds391
 PIN vss.gds392
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.866 2.9095 70.926 3.1095 ;
 END
 END vss.gds392
 PIN vss.gds393
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.034 2.9095 71.094 3.1095 ;
 END
 END vss.gds393
 PIN vss.gds394
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.202 2.9095 71.262 3.1095 ;
 END
 END vss.gds394
 PIN vss.gds395
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.538 2.9095 71.598 3.1095 ;
 END
 END vss.gds395
 PIN vss.gds396
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.706 2.9095 71.766 3.1095 ;
 END
 END vss.gds396
 PIN vss.gds397
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.874 2.9095 71.934 3.1095 ;
 END
 END vss.gds397
 PIN vss.gds398
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.21 2.9095 72.27 3.1095 ;
 END
 END vss.gds398
 PIN vss.gds399
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.378 2.9095 72.438 3.1095 ;
 END
 END vss.gds399
 PIN vss.gds400
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.546 2.9095 72.606 3.1095 ;
 END
 END vss.gds400
 PIN vss.gds401
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.882 2.9095 72.942 3.1095 ;
 END
 END vss.gds401
 PIN vss.gds402
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.05 2.9095 73.11 3.1095 ;
 END
 END vss.gds402
 PIN vss.gds403
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 2.9095 71.43 3.1095 ;
 END
 END vss.gds403
 PIN vss.gds404
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 2.9095 72.102 3.1095 ;
 END
 END vss.gds404
 PIN vss.gds405
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 2.9095 72.774 3.1095 ;
 END
 END vss.gds405
 PIN vss.gds406
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 2.9095 70.758 3.1095 ;
 END
 END vss.gds406
 PIN vss.gds407
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.554 2.9095 73.614 3.1095 ;
 END
 END vss.gds407
 PIN vss.gds408
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.722 2.9095 73.782 3.1095 ;
 END
 END vss.gds408
 PIN vss.gds409
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 2.9095 73.446 3.1095 ;
 END
 END vss.gds409
 PIN vss.gds410
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.218 2.9095 73.278 3.1095 ;
 END
 END vss.gds410
 PIN vss.gds411
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.89 2.9095 73.95 3.1095 ;
 END
 END vss.gds411
 PIN vss.gds412
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.394 2.9095 74.454 3.1095 ;
 END
 END vss.gds412
 PIN vss.gds413
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 2.9095 74.118 3.1095 ;
 END
 END vss.gds413
 PIN vss.gds414
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.562 2.9095 74.622 3.1095 ;
 END
 END vss.gds414
 PIN vss.gds415
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 2.9095 74.79 3.1095 ;
 END
 END vss.gds415
 PIN vss.gds416
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.226 2.9095 74.286 3.1095 ;
 END
 END vss.gds416
 PIN vss.gds417
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 5.953 2.962 6.153 ;
 END
 END vss.gds417
 PIN vss.gds418
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 7.213 2.962 7.413 ;
 END
 END vss.gds418
 PIN vss.gds419
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 7.437 0.942 7.637 ;
 END
 END vss.gds419
 PIN vss.gds420
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 9.332 3.142 9.532 ;
 END
 END vss.gds420
 PIN vss.gds421
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 9.733 2.962 9.933 ;
 END
 END vss.gds421
 PIN vss.gds422
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 8.473 2.962 8.673 ;
 END
 END vss.gds422
 PIN vss.gds423
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.286 7.843 3.326 8.043 ;
 END
 END vss.gds423
 PIN vss.gds424
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 7.843 4.194 8.043 ;
 END
 END vss.gds424
 PIN vss.gds425
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 7.843 5.074 8.043 ;
 END
 END vss.gds425
 PIN vss.gds426
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 7.5375 0.718 7.7375 ;
 END
 END vss.gds426
 PIN vss.gds427
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 5.552 3.142 5.752 ;
 END
 END vss.gds427
 PIN vss.gds428
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.442 7.437 4.482 7.637 ;
 END
 END vss.gds428
 PIN vss.gds429
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.57 7.64 4.61 7.84 ;
 END
 END vss.gds429
 PIN vss.gds430
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 7.437 4.882 7.637 ;
 END
 END vss.gds430
 PIN vss.gds431
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 7.638 0.602 7.838 ;
 END
 END vss.gds431
 PIN vss.gds432
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 8.072 3.142 8.272 ;
 END
 END vss.gds432
 PIN vss.gds433
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 7.8665 2.122 8.0665 ;
 END
 END vss.gds433
 PIN vss.gds434
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 7.981 1.282 8.181 ;
 END
 END vss.gds434
 PIN vss.gds435
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 8.2155 1.462 8.4155 ;
 END
 END vss.gds435
 PIN vss.gds436
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 6.812 3.142 7.012 ;
 END
 END vss.gds436
 PIN vss.gds437
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.414 8.119 3.454 8.319 ;
 END
 END vss.gds437
 PIN vss.gds438
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.562 8.119 3.602 8.319 ;
 END
 END vss.gds438
 PIN vss.gds439
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 7.778 2.302 7.978 ;
 END
 END vss.gds439
 PIN vss.gds440
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 7.7395 4.002 7.9395 ;
 END
 END vss.gds440
 PIN vss.gds441
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 7.7395 5.282 7.9395 ;
 END
 END vss.gds441
 PIN vss.gds442
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 7.824 0.29 8.024 ;
 END
 END vss.gds442
 PIN vss.gds443
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.754 7.843 3.794 8.043 ;
 END
 END vss.gds443
 PIN vss.gds444
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 2.408 5.9535 2.464 6.1535 ;
 RECT 2.576 5.9535 2.632 6.1535 ;
 RECT 2.996 5.9535 3.052 6.1535 ;
 RECT 3.332 6.045 3.388 6.245 ;
 RECT 3.5 6.0015 3.556 6.2015 ;
 RECT 0.98 5.8685 1.036 6.0685 ;
 RECT 2.072 5.869 2.128 6.069 ;
 RECT 2.576 7.2135 2.632 7.4135 ;
 RECT 2.408 7.2135 2.464 7.4135 ;
 RECT 2.996 7.2135 3.052 7.4135 ;
 RECT 3.332 7.305 3.388 7.505 ;
 RECT 2.576 8.4735 2.632 8.6735 ;
 RECT 2.408 8.4735 2.464 8.6735 ;
 RECT 2.996 8.4735 3.052 8.6735 ;
 RECT 3.332 8.565 3.388 8.765 ;
 RECT 2.408 9.7335 2.464 9.9335 ;
 RECT 2.576 9.7335 2.632 9.9335 ;
 RECT 2.996 9.7335 3.052 9.9335 ;
 RECT 3.332 9.825 3.388 10.025 ;
 RECT 3.5 9.7815 3.556 9.9815 ;
 RECT 0.98 9.6485 1.036 9.8485 ;
 RECT 2.072 9.649 2.128 9.849 ;
 RECT 0.812 8.565 0.868 8.765 ;
 RECT 3.5 7.2615 3.556 7.4615 ;
 RECT 0.98 7.1285 1.036 7.3285 ;
 RECT 2.072 7.129 2.128 7.329 ;
 RECT 0.392 7.219 0.448 7.419 ;
 RECT 0.812 7.305 0.868 7.505 ;
 RECT 0.644 7.219 0.7 7.419 ;
 RECT 1.232 7.219 1.288 7.419 ;
 RECT 1.4 7.219 1.456 7.419 ;
 RECT 1.568 7.219 1.624 7.419 ;
 RECT 1.82 7.219 1.876 7.419 ;
 RECT 2.24 7.219 2.296 7.419 ;
 RECT 2.744 7.129 2.8 7.329 ;
 RECT 3.164 7.219 3.22 7.419 ;
 RECT 3.5 8.5215 3.556 8.7215 ;
 RECT 0.392 8.479 0.448 8.679 ;
 RECT 0.644 8.479 0.7 8.679 ;
 RECT 1.232 8.479 1.288 8.679 ;
 RECT 0.98 8.3885 1.036 8.5885 ;
 RECT 1.4 8.479 1.456 8.679 ;
 RECT 1.568 8.479 1.624 8.679 ;
 RECT 2.072 8.389 2.128 8.589 ;
 RECT 1.82 8.479 1.876 8.679 ;
 RECT 2.744 8.389 2.8 8.589 ;
 RECT 3.164 8.479 3.22 8.679 ;
 RECT 2.24 8.479 2.296 8.679 ;
 RECT 0.392 9.739 0.448 9.939 ;
 RECT 0.812 9.825 0.868 10.025 ;
 RECT 0.644 9.739 0.7 9.939 ;
 RECT 1.232 9.739 1.288 9.939 ;
 RECT 1.4 9.739 1.456 9.939 ;
 RECT 1.568 9.739 1.624 9.939 ;
 RECT 1.82 9.739 1.876 9.939 ;
 RECT 2.24 9.739 2.296 9.939 ;
 RECT 2.744 9.649 2.8 9.849 ;
 RECT 3.164 9.739 3.22 9.939 ;
 RECT 3.92 9.739 3.976 9.939 ;
 RECT 3.752 10.009 3.808 10.209 ;
 RECT 4.508 9.9385 4.564 10.1385 ;
 RECT 3.92 8.479 3.976 8.679 ;
 RECT 3.752 8.749 3.808 8.949 ;
 RECT 4.508 8.6785 4.564 8.8785 ;
 RECT 3.92 7.219 3.976 7.419 ;
 RECT 3.752 7.489 3.808 7.689 ;
 RECT 4.508 7.4185 4.564 7.6185 ;
 RECT 0.392 5.959 0.448 6.159 ;
 RECT 0.812 6.045 0.868 6.245 ;
 RECT 0.644 5.959 0.7 6.159 ;
 RECT 1.232 5.959 1.288 6.159 ;
 RECT 1.4 5.959 1.456 6.159 ;
 RECT 1.568 5.959 1.624 6.159 ;
 RECT 1.82 5.959 1.876 6.159 ;
 RECT 2.24 5.959 2.296 6.159 ;
 RECT 2.744 5.869 2.8 6.069 ;
 RECT 3.164 5.959 3.22 6.159 ;
 RECT 3.92 5.959 3.976 6.159 ;
 RECT 3.752 6.229 3.808 6.429 ;
 RECT 4.508 6.1585 4.564 6.3585 ;
 END
 END vss.gds444
 PIN vss.gds445
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.134 8.0595 10.194 8.2595 ;
 END
 END vss.gds445
 PIN vss.gds446
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.966 8.0595 10.026 8.2595 ;
 END
 END vss.gds446
 PIN vss.gds447
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.798 8.0595 9.858 8.2595 ;
 END
 END vss.gds447
 PIN vss.gds448
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 8.0595 9.69 8.2595 ;
 END
 END vss.gds448
 PIN vss.gds449
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.462 8.0595 9.522 8.2595 ;
 END
 END vss.gds449
 PIN vss.gds450
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 8.0595 9.018 8.2595 ;
 END
 END vss.gds450
 PIN vss.gds451
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.79 8.0595 8.85 8.2595 ;
 END
 END vss.gds451
 PIN vss.gds452
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.622 8.0595 8.682 8.2595 ;
 END
 END vss.gds452
 PIN vss.gds453
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.454 8.0595 8.514 8.2595 ;
 END
 END vss.gds453
 PIN vss.gds454
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 7.843 5.474 8.043 ;
 END
 END vss.gds454
 PIN vss.gds455
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 8.0595 8.346 8.2595 ;
 END
 END vss.gds455
 PIN vss.gds456
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.118 8.0595 8.178 8.2595 ;
 END
 END vss.gds456
 PIN vss.gds457
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.95 8.0595 8.01 8.2595 ;
 END
 END vss.gds457
 PIN vss.gds458
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.294 8.0595 9.354 8.2595 ;
 END
 END vss.gds458
 PIN vss.gds459
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.782 8.0595 7.842 8.2595 ;
 END
 END vss.gds459
 PIN vss.gds460
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 8.0595 7.674 8.2595 ;
 END
 END vss.gds460
 PIN vss.gds461
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.126 8.0595 9.186 8.2595 ;
 END
 END vss.gds461
 PIN vss.gds462
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.446 8.0595 7.506 8.2595 ;
 END
 END vss.gds462
 PIN vss.gds463
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.278 8.0595 7.338 8.2595 ;
 END
 END vss.gds463
 PIN vss.gds464
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.11 8.0595 7.17 8.2595 ;
 END
 END vss.gds464
 PIN vss.gds465
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 7.843 5.73 8.043 ;
 END
 END vss.gds465
 PIN vss.gds466
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 7.843 5.986 8.043 ;
 END
 END vss.gds466
 PIN vss.gds467
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 7.639 6.434 7.839 ;
 END
 END vss.gds467
 PIN vss.gds468
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 7.64 6.178 7.84 ;
 END
 END vss.gds468
 PIN vss.gds469
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 6.608 10.009 6.664 10.209 ;
 RECT 6.524 9.732 6.58 9.932 ;
 RECT 6.692 9.882 6.748 10.082 ;
 RECT 6.692 8.622 6.748 8.822 ;
 RECT 6.524 8.472 6.58 8.672 ;
 RECT 6.608 8.749 6.664 8.949 ;
 RECT 6.692 7.362 6.748 7.562 ;
 RECT 6.524 7.212 6.58 7.412 ;
 RECT 6.608 7.489 6.664 7.689 ;
 RECT 6.608 6.229 6.664 6.429 ;
 RECT 6.524 5.952 6.58 6.152 ;
 RECT 6.692 6.102 6.748 6.302 ;
 END
 END vss.gds469
 PIN vss.gds470
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 7.758 14.87 7.958 ;
 END
 END vss.gds470
 PIN vss.gds471
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 6.458 13.898 6.658 ;
 END
 END vss.gds471
 PIN vss.gds472
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 6.498 14.87 6.698 ;
 END
 END vss.gds472
 PIN vss.gds473
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 8.978 13.898 9.178 ;
 END
 END vss.gds473
 PIN vss.gds474
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 9.018 14.87 9.218 ;
 END
 END vss.gds474
 PIN vss.gds475
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 10.238 13.898 10.438 ;
 END
 END vss.gds475
 PIN vss.gds476
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 10.278 14.87 10.478 ;
 END
 END vss.gds476
 PIN vss.gds477
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.15 8.0595 12.21 8.2595 ;
 END
 END vss.gds477
 PIN vss.gds478
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.982 8.0595 12.042 8.2595 ;
 END
 END vss.gds478
 PIN vss.gds479
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.814 8.0595 11.874 8.2595 ;
 END
 END vss.gds479
 PIN vss.gds480
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.478 8.0595 11.538 8.2595 ;
 END
 END vss.gds480
 PIN vss.gds481
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.31 8.0595 11.37 8.2595 ;
 END
 END vss.gds481
 PIN vss.gds482
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 8.1155 13.058 8.3155 ;
 END
 END vss.gds482
 PIN vss.gds483
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 8.0595 11.706 8.2595 ;
 END
 END vss.gds483
 PIN vss.gds484
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.142 8.0595 11.202 8.2595 ;
 END
 END vss.gds484
 PIN vss.gds485
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.806 8.0595 10.866 8.2595 ;
 END
 END vss.gds485
 PIN vss.gds486
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.638 8.0595 10.698 8.2595 ;
 END
 END vss.gds486
 PIN vss.gds487
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.47 8.0595 10.53 8.2595 ;
 END
 END vss.gds487
 PIN vss.gds488
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 8.0595 11.034 8.2595 ;
 END
 END vss.gds488
 PIN vss.gds489
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 8.0595 10.362 8.2595 ;
 END
 END vss.gds489
 PIN vss.gds490
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 8.1 15.162 8.3 ;
 END
 END vss.gds490
 PIN vss.gds491
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 8.1 14.498 8.3 ;
 END
 END vss.gds491
 PIN vss.gds492
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 7.718 13.898 7.918 ;
 END
 END vss.gds492
 PIN vss.gds493
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 8.0595 13.658 8.2595 ;
 END
 END vss.gds493
 PIN vss.gds494
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.262 8.112 13.318 8.312 ;
 END
 END vss.gds494
 PIN vss.gds495
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 7.981 12.378 8.181 ;
 END
 END vss.gds495
 PIN vss.gds496
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 7.843 12.59 8.043 ;
 END
 END vss.gds496
 PIN vss.gds497
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 7.9635 12.818 8.1635 ;
 END
 END vss.gds497
 PIN vss.gds498
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 14 9.156 14.056 9.329 ;
 RECT 14.168 9.129 14.224 9.329 ;
 RECT 14 6.636 14.056 6.809 ;
 RECT 14.168 6.609 14.224 6.809 ;
 RECT 14 7.896 14.056 8.069 ;
 RECT 14.168 7.869 14.224 8.069 ;
 RECT 14 10.416 14.056 10.589 ;
 RECT 14.168 10.389 14.224 10.589 ;
 RECT 14.336 5.969 14.392 6.169 ;
 RECT 14.168 5.969 14.224 6.169 ;
 RECT 14.336 8.489 14.392 8.689 ;
 RECT 14.168 8.489 14.224 8.689 ;
 RECT 14.336 9.749 14.392 9.949 ;
 RECT 14.168 9.749 14.224 9.949 ;
 RECT 13.664 9.883 13.72 10.083 ;
 RECT 15.008 9.959 15.064 10.159 ;
 RECT 14.84 10.433 14.896 10.598 ;
 RECT 14.672 10.433 14.728 10.598 ;
 RECT 14.336 7.229 14.392 7.429 ;
 RECT 14.168 7.229 14.224 7.429 ;
 RECT 15.008 7.439 15.064 7.639 ;
 RECT 14.84 7.913 14.896 8.078 ;
 RECT 14.672 7.913 14.728 8.078 ;
 RECT 15.008 6.179 15.064 6.379 ;
 RECT 14.84 6.653 14.896 6.818 ;
 RECT 14.672 6.653 14.728 6.818 ;
 RECT 13.664 6.103 13.72 6.303 ;
 RECT 13.664 8.623 13.72 8.823 ;
 RECT 15.008 8.699 15.064 8.899 ;
 RECT 14.84 9.173 14.896 9.338 ;
 RECT 14.672 9.173 14.728 9.338 ;
 RECT 13.664 7.363 13.72 7.563 ;
 RECT 15.176 8.1395 15.232 8.3395 ;
 RECT 12.824 7.924 12.88 8.124 ;
 RECT 13.496 7.935 13.552 8.135 ;
 RECT 12.488 7.954 12.544 8.154 ;
 RECT 13.328 7.873 13.384 8.073 ;
 RECT 13.16 7.924 13.216 8.124 ;
 RECT 12.992 7.924 13.048 8.124 ;
 RECT 12.656 7.954 12.712 8.154 ;
 END
 END vss.gds498
 PIN vss.gds499
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 7.956 15.418 8.156 ;
 END
 END vss.gds499
 PIN vss.gds500
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 8.0595 20.274 8.2595 ;
 END
 END vss.gds500
 PIN vss.gds501
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 8.0595 18.93 8.2595 ;
 END
 END vss.gds501
 PIN vss.gds502
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.038 8.0595 19.098 8.2595 ;
 END
 END vss.gds502
 PIN vss.gds503
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.206 8.0595 19.266 8.2595 ;
 END
 END vss.gds503
 PIN vss.gds504
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.374 8.0595 19.434 8.2595 ;
 END
 END vss.gds504
 PIN vss.gds505
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 8.0595 19.602 8.2595 ;
 END
 END vss.gds505
 PIN vss.gds506
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 7.9635 17.314 8.1635 ;
 END
 END vss.gds506
 PIN vss.gds507
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 8.0185 16.994 8.2185 ;
 END
 END vss.gds507
 PIN vss.gds508
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.71 8.0595 19.77 8.2595 ;
 END
 END vss.gds508
 PIN vss.gds509
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.878 8.0595 19.938 8.2595 ;
 END
 END vss.gds509
 PIN vss.gds510
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 9.733 16.146 9.933 ;
 END
 END vss.gds510
 PIN vss.gds511
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 7.213 16.146 7.413 ;
 END
 END vss.gds511
 PIN vss.gds512
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 8.473 16.146 8.673 ;
 END
 END vss.gds512
 PIN vss.gds513
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 5.953 16.146 6.153 ;
 END
 END vss.gds513
 PIN vss.gds514
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 8.1 15.842 8.3 ;
 END
 END vss.gds514
 PIN vss.gds515
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 8.112 16.814 8.312 ;
 END
 END vss.gds515
 PIN vss.gds516
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.046 8.0595 20.106 8.2595 ;
 END
 END vss.gds516
 PIN vss.gds517
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.702 8.0595 18.762 8.2595 ;
 END
 END vss.gds517
 PIN vss.gds518
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.534 8.0595 18.594 8.2595 ;
 END
 END vss.gds518
 PIN vss.gds519
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.366 8.0595 18.426 8.2595 ;
 END
 END vss.gds519
 PIN vss.gds520
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 7.981 18.258 8.181 ;
 END
 END vss.gds520
 PIN vss.gds521
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 7.9635 17.834 8.1635 ;
 END
 END vss.gds521
 PIN vss.gds522
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.438 8.1155 17.494 8.3155 ;
 END
 END vss.gds522
 PIN vss.gds523
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 7.8665 16.49 8.0665 ;
 END
 END vss.gds523
 PIN vss.gds524
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.986 7.843 18.026 8.043 ;
 END
 END vss.gds524
 PIN vss.gds525
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 15.596 6.88 15.652 7.08 ;
 RECT 15.848 6.883 15.904 7.083 ;
 RECT 15.596 8.14 15.652 8.34 ;
 RECT 15.848 8.143 15.904 8.343 ;
 RECT 16.52 9.176 16.576 9.329 ;
 RECT 15.764 9.173 15.82 9.338 ;
 RECT 15.596 9.173 15.652 9.338 ;
 RECT 15.596 5.62 15.652 5.82 ;
 RECT 15.848 5.623 15.904 5.823 ;
 RECT 16.52 6.656 16.576 6.809 ;
 RECT 15.764 6.653 15.82 6.818 ;
 RECT 15.596 6.653 15.652 6.818 ;
 RECT 16.52 7.916 16.576 8.069 ;
 RECT 15.764 7.913 15.82 8.078 ;
 RECT 15.596 7.913 15.652 8.078 ;
 RECT 15.596 9.4 15.652 9.6 ;
 RECT 15.848 9.403 15.904 9.603 ;
 RECT 16.52 10.436 16.576 10.589 ;
 RECT 15.764 10.433 15.82 10.598 ;
 RECT 15.596 10.433 15.652 10.598 ;
 RECT 16.352 10.0595 16.408 10.2595 ;
 RECT 16.856 9.8075 16.912 10.0075 ;
 RECT 16.352 8.7995 16.408 8.9995 ;
 RECT 16.856 8.5475 16.912 8.7475 ;
 RECT 15.428 9.959 15.484 10.159 ;
 RECT 15.428 7.439 15.484 7.639 ;
 RECT 15.428 6.179 15.484 6.379 ;
 RECT 16.352 6.2795 16.408 6.4795 ;
 RECT 16.856 6.0275 16.912 6.2275 ;
 RECT 15.428 8.699 15.484 8.899 ;
 RECT 16.352 7.5395 16.408 7.7395 ;
 RECT 16.856 7.2875 16.912 7.4875 ;
 RECT 17.864 7.954 17.92 8.154 ;
 RECT 17.696 7.9615 17.752 8.1615 ;
 RECT 17.528 7.954 17.584 8.154 ;
 RECT 17.36 7.954 17.416 8.154 ;
 RECT 17.192 7.954 17.248 8.154 ;
 RECT 18.032 7.954 18.088 8.154 ;
 RECT 17.024 8.069 17.08 8.269 ;
 END
 END vss.gds525
 PIN vss.gds526
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.17 8.0595 25.23 8.2595 ;
 END
 END vss.gds526
 PIN vss.gds527
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.002 8.0595 25.062 8.2595 ;
 END
 END vss.gds527
 PIN vss.gds528
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.834 8.0595 24.894 8.2595 ;
 END
 END vss.gds528
 PIN vss.gds529
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.498 8.0595 24.558 8.2595 ;
 END
 END vss.gds529
 PIN vss.gds530
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.33 8.0595 24.39 8.2595 ;
 END
 END vss.gds530
 PIN vss.gds531
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.162 8.0595 24.222 8.2595 ;
 END
 END vss.gds531
 PIN vss.gds532
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.382 8.0595 20.442 8.2595 ;
 END
 END vss.gds532
 PIN vss.gds533
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.55 8.0595 20.61 8.2595 ;
 END
 END vss.gds533
 PIN vss.gds534
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.718 8.0595 20.778 8.2595 ;
 END
 END vss.gds534
 PIN vss.gds535
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.054 8.0595 21.114 8.2595 ;
 END
 END vss.gds535
 PIN vss.gds536
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.222 8.0595 21.282 8.2595 ;
 END
 END vss.gds536
 PIN vss.gds537
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.39 8.0595 21.45 8.2595 ;
 END
 END vss.gds537
 PIN vss.gds538
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.726 8.0595 21.786 8.2595 ;
 END
 END vss.gds538
 PIN vss.gds539
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.894 8.0595 21.954 8.2595 ;
 END
 END vss.gds539
 PIN vss.gds540
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.062 8.0595 22.122 8.2595 ;
 END
 END vss.gds540
 PIN vss.gds541
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.398 8.0595 22.458 8.2595 ;
 END
 END vss.gds541
 PIN vss.gds542
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.566 8.0595 22.626 8.2595 ;
 END
 END vss.gds542
 PIN vss.gds543
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.734 8.0595 22.794 8.2595 ;
 END
 END vss.gds543
 PIN vss.gds544
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 8.0595 24.726 8.2595 ;
 END
 END vss.gds544
 PIN vss.gds545
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 8.0595 21.618 8.2595 ;
 END
 END vss.gds545
 PIN vss.gds546
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 8.0595 20.946 8.2595 ;
 END
 END vss.gds546
 PIN vss.gds547
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 8.0595 22.29 8.2595 ;
 END
 END vss.gds547
 PIN vss.gds548
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 8.0595 22.962 8.2595 ;
 END
 END vss.gds548
 PIN vss.gds549
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.07 8.0595 23.13 8.2595 ;
 END
 END vss.gds549
 PIN vss.gds550
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.238 8.0595 23.298 8.2595 ;
 END
 END vss.gds550
 PIN vss.gds551
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.406 8.0595 23.466 8.2595 ;
 END
 END vss.gds551
 PIN vss.gds552
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 8.0595 23.634 8.2595 ;
 END
 END vss.gds552
 PIN vss.gds553
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 23.912 9.896 23.968 10.096 ;
 RECT 23.912 8.636 23.968 8.836 ;
 RECT 23.912 7.376 23.968 7.576 ;
 RECT 23.912 6.116 23.968 6.316 ;
 RECT 23.744 8.006 23.8 8.206 ;
 END
 END vss.gds553
 PIN vss.gds554
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.202 8.0595 29.262 8.2595 ;
 END
 END vss.gds554
 PIN vss.gds555
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.034 8.0595 29.094 8.2595 ;
 END
 END vss.gds555
 PIN vss.gds556
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.866 8.0595 28.926 8.2595 ;
 END
 END vss.gds556
 PIN vss.gds557
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.53 8.0595 28.59 8.2595 ;
 END
 END vss.gds557
 PIN vss.gds558
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.362 8.0595 28.422 8.2595 ;
 END
 END vss.gds558
 PIN vss.gds559
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.194 8.0595 28.254 8.2595 ;
 END
 END vss.gds559
 PIN vss.gds560
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.858 8.0595 27.918 8.2595 ;
 END
 END vss.gds560
 PIN vss.gds561
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.69 8.0595 27.75 8.2595 ;
 END
 END vss.gds561
 PIN vss.gds562
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.522 8.0595 27.582 8.2595 ;
 END
 END vss.gds562
 PIN vss.gds563
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.186 8.0595 27.246 8.2595 ;
 END
 END vss.gds563
 PIN vss.gds564
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.018 8.0595 27.078 8.2595 ;
 END
 END vss.gds564
 PIN vss.gds565
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.85 8.0595 26.91 8.2595 ;
 END
 END vss.gds565
 PIN vss.gds566
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.514 8.0595 26.574 8.2595 ;
 END
 END vss.gds566
 PIN vss.gds567
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.346 8.0595 26.406 8.2595 ;
 END
 END vss.gds567
 PIN vss.gds568
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.178 8.0595 26.238 8.2595 ;
 END
 END vss.gds568
 PIN vss.gds569
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.842 8.0595 25.902 8.2595 ;
 END
 END vss.gds569
 PIN vss.gds570
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.674 8.0595 25.734 8.2595 ;
 END
 END vss.gds570
 PIN vss.gds571
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.506 8.0595 25.566 8.2595 ;
 END
 END vss.gds571
 PIN vss.gds572
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 8.0595 28.758 8.2595 ;
 END
 END vss.gds572
 PIN vss.gds573
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 8.0595 28.086 8.2595 ;
 END
 END vss.gds573
 PIN vss.gds574
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 8.0595 27.414 8.2595 ;
 END
 END vss.gds574
 PIN vss.gds575
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 8.0595 26.742 8.2595 ;
 END
 END vss.gds575
 PIN vss.gds576
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 8.0595 26.07 8.2595 ;
 END
 END vss.gds576
 PIN vss.gds577
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 8.0595 25.398 8.2595 ;
 END
 END vss.gds577
 PIN vss.gds578
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 7.981 29.43 8.181 ;
 END
 END vss.gds578
 PIN vss.gds579
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 8.1155 30.11 8.3155 ;
 END
 END vss.gds579
 PIN vss.gds580
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 7.9635 29.87 8.1635 ;
 END
 END vss.gds580
 PIN vss.gds581
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 7.843 29.642 8.043 ;
 END
 END vss.gds581
 PIN vss.gds582
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.876 7.924 29.932 8.124 ;
 RECT 30.212 7.924 30.268 8.124 ;
 RECT 29.54 7.954 29.596 8.154 ;
 RECT 30.044 7.924 30.1 8.124 ;
 RECT 29.708 7.954 29.764 8.154 ;
 END
 END vss.gds582
 PIN vss.gds583
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 7.758 31.922 7.958 ;
 END
 END vss.gds583
 PIN vss.gds584
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 7.718 30.95 7.918 ;
 END
 END vss.gds584
 PIN vss.gds585
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 6.498 31.922 6.698 ;
 END
 END vss.gds585
 PIN vss.gds586
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 8.978 30.95 9.178 ;
 END
 END vss.gds586
 PIN vss.gds587
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 9.018 31.922 9.218 ;
 END
 END vss.gds587
 PIN vss.gds588
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 10.238 30.95 10.438 ;
 END
 END vss.gds588
 PIN vss.gds589
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 10.278 31.922 10.478 ;
 END
 END vss.gds589
 PIN vss.gds590
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.314 8.112 30.37 8.312 ;
 END
 END vss.gds590
 PIN vss.gds591
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 8.1 32.214 8.3 ;
 END
 END vss.gds591
 PIN vss.gds592
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 8.0185 34.046 8.2185 ;
 END
 END vss.gds592
 PIN vss.gds593
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 8.0595 30.71 8.2595 ;
 END
 END vss.gds593
 PIN vss.gds594
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 8.1 32.894 8.3 ;
 END
 END vss.gds594
 PIN vss.gds595
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 9.733 33.198 9.933 ;
 END
 END vss.gds595
 PIN vss.gds596
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 8.473 33.198 8.673 ;
 END
 END vss.gds596
 PIN vss.gds597
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 7.8665 33.542 8.0665 ;
 END
 END vss.gds597
 PIN vss.gds598
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 8.1 31.55 8.3 ;
 END
 END vss.gds598
 PIN vss.gds599
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 8.112 33.866 8.312 ;
 END
 END vss.gds599
 PIN vss.gds600
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 5.953 33.198 6.153 ;
 END
 END vss.gds600
 PIN vss.gds601
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 7.213 33.198 7.413 ;
 END
 END vss.gds601
 PIN vss.gds602
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 7.9635 34.886 8.1635 ;
 END
 END vss.gds602
 PIN vss.gds603
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.49 8.1155 34.546 8.3155 ;
 END
 END vss.gds603
 PIN vss.gds604
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 7.956 32.47 8.156 ;
 END
 END vss.gds604
 PIN vss.gds605
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 6.458 30.95 6.658 ;
 END
 END vss.gds605
 PIN vss.gds606
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 7.9635 34.366 8.1635 ;
 END
 END vss.gds606
 PIN vss.gds607
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.038 7.843 35.078 8.043 ;
 END
 END vss.gds607
 PIN vss.gds608
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 32.648 6.88 32.704 7.08 ;
 RECT 32.9 6.883 32.956 7.083 ;
 RECT 33.572 9.176 33.628 9.329 ;
 RECT 31.052 9.156 31.108 9.329 ;
 RECT 31.22 9.129 31.276 9.329 ;
 RECT 32.816 9.173 32.872 9.338 ;
 RECT 32.648 9.173 32.704 9.338 ;
 RECT 31.892 9.173 31.948 9.338 ;
 RECT 31.724 9.173 31.78 9.338 ;
 RECT 32.648 5.62 32.704 5.82 ;
 RECT 32.9 5.623 32.956 5.823 ;
 RECT 33.572 6.656 33.628 6.809 ;
 RECT 31.052 6.636 31.108 6.809 ;
 RECT 31.22 6.609 31.276 6.809 ;
 RECT 32.816 6.653 32.872 6.818 ;
 RECT 32.648 6.653 32.704 6.818 ;
 RECT 31.892 6.653 31.948 6.818 ;
 RECT 31.724 6.653 31.78 6.818 ;
 RECT 33.572 7.916 33.628 8.069 ;
 RECT 31.052 7.896 31.108 8.069 ;
 RECT 31.22 7.869 31.276 8.069 ;
 RECT 32.816 7.913 32.872 8.078 ;
 RECT 32.648 7.913 32.704 8.078 ;
 RECT 31.892 7.913 31.948 8.078 ;
 RECT 31.724 7.913 31.78 8.078 ;
 RECT 33.572 10.436 33.628 10.589 ;
 RECT 31.052 10.416 31.108 10.589 ;
 RECT 31.22 10.389 31.276 10.589 ;
 RECT 32.816 10.433 32.872 10.598 ;
 RECT 32.648 10.433 32.704 10.598 ;
 RECT 31.892 10.433 31.948 10.598 ;
 RECT 31.724 10.433 31.78 10.598 ;
 RECT 32.648 8.14 32.704 8.34 ;
 RECT 32.9 8.143 32.956 8.343 ;
 RECT 32.648 9.4 32.704 9.6 ;
 RECT 32.9 9.403 32.956 9.603 ;
 RECT 31.388 8.489 31.444 8.689 ;
 RECT 31.22 8.489 31.276 8.689 ;
 RECT 33.404 8.7995 33.46 8.9995 ;
 RECT 33.908 8.5475 33.964 8.7475 ;
 RECT 33.908 9.8075 33.964 10.0075 ;
 RECT 33.404 10.0595 33.46 10.2595 ;
 RECT 32.06 9.959 32.116 10.159 ;
 RECT 32.48 9.959 32.536 10.159 ;
 RECT 31.388 9.749 31.444 9.949 ;
 RECT 31.22 9.749 31.276 9.949 ;
 RECT 30.716 9.883 30.772 10.083 ;
 RECT 31.388 5.969 31.444 6.169 ;
 RECT 31.22 5.969 31.276 6.169 ;
 RECT 32.06 6.179 32.116 6.379 ;
 RECT 32.48 6.179 32.536 6.379 ;
 RECT 33.908 7.2875 33.964 7.4875 ;
 RECT 33.404 7.5395 33.46 7.7395 ;
 RECT 32.06 7.439 32.116 7.639 ;
 RECT 32.48 7.439 32.536 7.639 ;
 RECT 31.388 7.229 31.444 7.429 ;
 RECT 31.22 7.229 31.276 7.429 ;
 RECT 30.716 7.363 30.772 7.563 ;
 RECT 30.716 8.623 30.772 8.823 ;
 RECT 32.06 8.699 32.116 8.899 ;
 RECT 32.48 8.699 32.536 8.899 ;
 RECT 30.716 6.103 30.772 6.303 ;
 RECT 33.404 6.2795 33.46 6.4795 ;
 RECT 33.908 6.0275 33.964 6.2275 ;
 RECT 30.548 7.935 30.604 8.135 ;
 RECT 30.38 7.873 30.436 8.073 ;
 RECT 32.228 8.1395 32.284 8.3395 ;
 RECT 34.916 7.954 34.972 8.154 ;
 RECT 34.748 7.9615 34.804 8.1615 ;
 RECT 34.58 7.954 34.636 8.154 ;
 RECT 34.412 7.954 34.468 8.154 ;
 RECT 34.244 7.954 34.3 8.154 ;
 RECT 35.084 7.954 35.14 8.154 ;
 RECT 34.076 8.069 34.132 8.269 ;
 END
 END vss.gds608
 PIN vss.gds609
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.122 8.0595 40.182 8.2595 ;
 END
 END vss.gds609
 PIN vss.gds610
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.754 8.0595 35.814 8.2595 ;
 END
 END vss.gds610
 PIN vss.gds611
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.09 8.0595 36.15 8.2595 ;
 END
 END vss.gds611
 PIN vss.gds612
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.258 8.0595 36.318 8.2595 ;
 END
 END vss.gds612
 PIN vss.gds613
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.426 8.0595 36.486 8.2595 ;
 END
 END vss.gds613
 PIN vss.gds614
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.762 8.0595 36.822 8.2595 ;
 END
 END vss.gds614
 PIN vss.gds615
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.93 8.0595 36.99 8.2595 ;
 END
 END vss.gds615
 PIN vss.gds616
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.098 8.0595 37.158 8.2595 ;
 END
 END vss.gds616
 PIN vss.gds617
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.434 8.0595 37.494 8.2595 ;
 END
 END vss.gds617
 PIN vss.gds618
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.602 8.0595 37.662 8.2595 ;
 END
 END vss.gds618
 PIN vss.gds619
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.77 8.0595 37.83 8.2595 ;
 END
 END vss.gds619
 PIN vss.gds620
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.106 8.0595 38.166 8.2595 ;
 END
 END vss.gds620
 PIN vss.gds621
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.274 8.0595 38.334 8.2595 ;
 END
 END vss.gds621
 PIN vss.gds622
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 8.0595 36.654 8.2595 ;
 END
 END vss.gds622
 PIN vss.gds623
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 8.0595 37.326 8.2595 ;
 END
 END vss.gds623
 PIN vss.gds624
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 8.0595 37.998 8.2595 ;
 END
 END vss.gds624
 PIN vss.gds625
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.442 8.0595 38.502 8.2595 ;
 END
 END vss.gds625
 PIN vss.gds626
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 8.0595 38.67 8.2595 ;
 END
 END vss.gds626
 PIN vss.gds627
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.778 8.0595 38.838 8.2595 ;
 END
 END vss.gds627
 PIN vss.gds628
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 8.0595 35.982 8.2595 ;
 END
 END vss.gds628
 PIN vss.gds629
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.946 8.0595 39.006 8.2595 ;
 END
 END vss.gds629
 PIN vss.gds630
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.586 8.0595 35.646 8.2595 ;
 END
 END vss.gds630
 PIN vss.gds631
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.45 8.0595 39.51 8.2595 ;
 END
 END vss.gds631
 PIN vss.gds632
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.618 8.0595 39.678 8.2595 ;
 END
 END vss.gds632
 PIN vss.gds633
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.114 8.0595 39.174 8.2595 ;
 END
 END vss.gds633
 PIN vss.gds634
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.786 8.0595 39.846 8.2595 ;
 END
 END vss.gds634
 PIN vss.gds635
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 8.0595 40.014 8.2595 ;
 END
 END vss.gds635
 PIN vss.gds636
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.418 8.0595 35.478 8.2595 ;
 END
 END vss.gds636
 PIN vss.gds637
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 7.981 35.31 8.181 ;
 END
 END vss.gds637
 PIN vss.gds638
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 8.0595 39.342 8.2595 ;
 END
 END vss.gds638
 PIN vss.gds639
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.91 8.0595 44.97 8.2595 ;
 END
 END vss.gds639
 PIN vss.gds640
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.742 8.0595 44.802 8.2595 ;
 END
 END vss.gds640
 PIN vss.gds641
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.574 8.0595 44.634 8.2595 ;
 END
 END vss.gds641
 PIN vss.gds642
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.238 8.0595 44.298 8.2595 ;
 END
 END vss.gds642
 PIN vss.gds643
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.07 8.0595 44.13 8.2595 ;
 END
 END vss.gds643
 PIN vss.gds644
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.902 8.0595 43.962 8.2595 ;
 END
 END vss.gds644
 PIN vss.gds645
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.566 8.0595 43.626 8.2595 ;
 END
 END vss.gds645
 PIN vss.gds646
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.398 8.0595 43.458 8.2595 ;
 END
 END vss.gds646
 PIN vss.gds647
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.23 8.0595 43.29 8.2595 ;
 END
 END vss.gds647
 PIN vss.gds648
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.894 8.0595 42.954 8.2595 ;
 END
 END vss.gds648
 PIN vss.gds649
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.726 8.0595 42.786 8.2595 ;
 END
 END vss.gds649
 PIN vss.gds650
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.558 8.0595 42.618 8.2595 ;
 END
 END vss.gds650
 PIN vss.gds651
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.222 8.0595 42.282 8.2595 ;
 END
 END vss.gds651
 PIN vss.gds652
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.054 8.0595 42.114 8.2595 ;
 END
 END vss.gds652
 PIN vss.gds653
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.886 8.0595 41.946 8.2595 ;
 END
 END vss.gds653
 PIN vss.gds654
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.55 8.0595 41.61 8.2595 ;
 END
 END vss.gds654
 PIN vss.gds655
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.382 8.0595 41.442 8.2595 ;
 END
 END vss.gds655
 PIN vss.gds656
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.214 8.0595 41.274 8.2595 ;
 END
 END vss.gds656
 PIN vss.gds657
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.29 8.0595 40.35 8.2595 ;
 END
 END vss.gds657
 PIN vss.gds658
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.458 8.0595 40.518 8.2595 ;
 END
 END vss.gds658
 PIN vss.gds659
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 8.0595 45.138 8.2595 ;
 END
 END vss.gds659
 PIN vss.gds660
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 8.0595 44.466 8.2595 ;
 END
 END vss.gds660
 PIN vss.gds661
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 8.0595 43.794 8.2595 ;
 END
 END vss.gds661
 PIN vss.gds662
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 8.0595 43.122 8.2595 ;
 END
 END vss.gds662
 PIN vss.gds663
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 8.0595 42.45 8.2595 ;
 END
 END vss.gds663
 PIN vss.gds664
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 8.0595 41.778 8.2595 ;
 END
 END vss.gds664
 PIN vss.gds665
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 8.0595 40.686 8.2595 ;
 END
 END vss.gds665
 PIN vss.gds666
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 40.964 8.636 41.02 8.836 ;
 RECT 40.964 9.896 41.02 10.096 ;
 RECT 40.964 6.116 41.02 6.316 ;
 RECT 40.964 7.376 41.02 7.576 ;
 RECT 40.796 8.006 40.852 8.206 ;
 END
 END vss.gds666
 PIN vss.gds667
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 7.758 48.974 7.958 ;
 END
 END vss.gds667
 PIN vss.gds668
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 6.498 48.974 6.698 ;
 END
 END vss.gds668
 PIN vss.gds669
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 9.018 48.974 9.218 ;
 END
 END vss.gds669
 PIN vss.gds670
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 6.458 48.002 6.658 ;
 END
 END vss.gds670
 PIN vss.gds671
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 10.278 48.974 10.478 ;
 END
 END vss.gds671
 PIN vss.gds672
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 8.978 48.002 9.178 ;
 END
 END vss.gds672
 PIN vss.gds673
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 10.238 48.002 10.438 ;
 END
 END vss.gds673
 PIN vss.gds674
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.366 8.112 47.422 8.312 ;
 END
 END vss.gds674
 PIN vss.gds675
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.254 8.0595 46.314 8.2595 ;
 END
 END vss.gds675
 PIN vss.gds676
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.086 8.0595 46.146 8.2595 ;
 END
 END vss.gds676
 PIN vss.gds677
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.918 8.0595 45.978 8.2595 ;
 END
 END vss.gds677
 PIN vss.gds678
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.582 8.0595 45.642 8.2595 ;
 END
 END vss.gds678
 PIN vss.gds679
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.414 8.0595 45.474 8.2595 ;
 END
 END vss.gds679
 PIN vss.gds680
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.246 8.0595 45.306 8.2595 ;
 END
 END vss.gds680
 PIN vss.gds681
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 8.1155 47.162 8.3155 ;
 END
 END vss.gds681
 PIN vss.gds682
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 7.981 46.482 8.181 ;
 END
 END vss.gds682
 PIN vss.gds683
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 8.0595 45.81 8.2595 ;
 END
 END vss.gds683
 PIN vss.gds684
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 7.9635 46.922 8.1635 ;
 END
 END vss.gds684
 PIN vss.gds685
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 7.843 46.694 8.043 ;
 END
 END vss.gds685
 PIN vss.gds686
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 8.0595 47.762 8.2595 ;
 END
 END vss.gds686
 PIN vss.gds687
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 8.1 49.266 8.3 ;
 END
 END vss.gds687
 PIN vss.gds688
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 8.1 48.602 8.3 ;
 END
 END vss.gds688
 PIN vss.gds689
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 8.1 49.946 8.3 ;
 END
 END vss.gds689
 PIN vss.gds690
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 9.733 50.25 9.933 ;
 END
 END vss.gds690
 PIN vss.gds691
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 8.473 50.25 8.673 ;
 END
 END vss.gds691
 PIN vss.gds692
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 7.213 50.25 7.413 ;
 END
 END vss.gds692
 PIN vss.gds693
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 5.953 50.25 6.153 ;
 END
 END vss.gds693
 PIN vss.gds694
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 7.718 48.002 7.918 ;
 END
 END vss.gds694
 PIN vss.gds695
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 7.956 49.522 8.156 ;
 END
 END vss.gds695
 PIN vss.gds696
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 48.104 9.156 48.16 9.329 ;
 RECT 48.272 9.129 48.328 9.329 ;
 RECT 49.868 9.173 49.924 9.338 ;
 RECT 49.7 9.173 49.756 9.338 ;
 RECT 48.944 9.173 49 9.338 ;
 RECT 48.776 9.173 48.832 9.338 ;
 RECT 48.104 6.636 48.16 6.809 ;
 RECT 48.272 6.609 48.328 6.809 ;
 RECT 49.868 6.653 49.924 6.818 ;
 RECT 49.7 6.653 49.756 6.818 ;
 RECT 48.944 6.653 49 6.818 ;
 RECT 48.776 6.653 48.832 6.818 ;
 RECT 48.104 7.896 48.16 8.069 ;
 RECT 48.272 7.869 48.328 8.069 ;
 RECT 49.868 7.913 49.924 8.078 ;
 RECT 49.7 7.913 49.756 8.078 ;
 RECT 48.944 7.913 49 8.078 ;
 RECT 48.776 7.913 48.832 8.078 ;
 RECT 48.104 10.416 48.16 10.589 ;
 RECT 48.272 10.389 48.328 10.589 ;
 RECT 49.868 10.433 49.924 10.598 ;
 RECT 49.7 10.433 49.756 10.598 ;
 RECT 48.944 10.433 49 10.598 ;
 RECT 48.776 10.433 48.832 10.598 ;
 RECT 49.7 5.62 49.756 5.82 ;
 RECT 49.952 5.623 50.008 5.823 ;
 RECT 49.7 6.88 49.756 7.08 ;
 RECT 49.952 6.883 50.008 7.083 ;
 RECT 49.7 9.4 49.756 9.6 ;
 RECT 49.952 9.403 50.008 9.603 ;
 RECT 49.7 8.14 49.756 8.34 ;
 RECT 49.952 8.143 50.008 8.343 ;
 RECT 48.44 9.749 48.496 9.949 ;
 RECT 48.272 9.749 48.328 9.949 ;
 RECT 47.768 9.883 47.824 10.083 ;
 RECT 49.112 9.959 49.168 10.159 ;
 RECT 49.532 9.959 49.588 10.159 ;
 RECT 48.44 7.229 48.496 7.429 ;
 RECT 48.272 7.229 48.328 7.429 ;
 RECT 49.112 7.439 49.168 7.639 ;
 RECT 49.532 7.439 49.588 7.639 ;
 RECT 48.44 8.489 48.496 8.689 ;
 RECT 48.272 8.489 48.328 8.689 ;
 RECT 47.768 8.623 47.824 8.823 ;
 RECT 49.112 8.699 49.168 8.899 ;
 RECT 49.532 8.699 49.588 8.899 ;
 RECT 47.768 7.363 47.824 7.563 ;
 RECT 49.112 6.179 49.168 6.379 ;
 RECT 49.532 6.179 49.588 6.379 ;
 RECT 48.44 5.969 48.496 6.169 ;
 RECT 48.272 5.969 48.328 6.169 ;
 RECT 47.768 6.103 47.824 6.303 ;
 RECT 47.6 7.935 47.656 8.135 ;
 RECT 47.432 7.873 47.488 8.073 ;
 RECT 47.264 7.924 47.32 8.124 ;
 RECT 46.928 7.924 46.984 8.124 ;
 RECT 47.096 7.924 47.152 8.124 ;
 RECT 49.28 8.1395 49.336 8.3395 ;
 RECT 46.592 7.954 46.648 8.154 ;
 RECT 46.76 7.954 46.816 8.154 ;
 END
 END vss.gds696
 PIN vss.gds697
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.638 8.0595 52.698 8.2595 ;
 END
 END vss.gds697
 PIN vss.gds698
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.806 8.0595 52.866 8.2595 ;
 END
 END vss.gds698
 PIN vss.gds699
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.142 8.0595 53.202 8.2595 ;
 END
 END vss.gds699
 PIN vss.gds700
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.31 8.0595 53.37 8.2595 ;
 END
 END vss.gds700
 PIN vss.gds701
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.478 8.0595 53.538 8.2595 ;
 END
 END vss.gds701
 PIN vss.gds702
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.814 8.0595 53.874 8.2595 ;
 END
 END vss.gds702
 PIN vss.gds703
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.982 8.0595 54.042 8.2595 ;
 END
 END vss.gds703
 PIN vss.gds704
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.15 8.0595 54.21 8.2595 ;
 END
 END vss.gds704
 PIN vss.gds705
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.486 8.0595 54.546 8.2595 ;
 END
 END vss.gds705
 PIN vss.gds706
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.654 8.0595 54.714 8.2595 ;
 END
 END vss.gds706
 PIN vss.gds707
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.822 8.0595 54.882 8.2595 ;
 END
 END vss.gds707
 PIN vss.gds708
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.158 8.0595 55.218 8.2595 ;
 END
 END vss.gds708
 PIN vss.gds709
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 8.0595 55.05 8.2595 ;
 END
 END vss.gds709
 PIN vss.gds710
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 8.0595 54.378 8.2595 ;
 END
 END vss.gds710
 PIN vss.gds711
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 8.112 50.918 8.312 ;
 END
 END vss.gds711
 PIN vss.gds712
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 8.0595 53.706 8.2595 ;
 END
 END vss.gds712
 PIN vss.gds713
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 8.0185 51.098 8.2185 ;
 END
 END vss.gds713
 PIN vss.gds714
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 8.0595 53.034 8.2595 ;
 END
 END vss.gds714
 PIN vss.gds715
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 7.9635 51.938 8.1635 ;
 END
 END vss.gds715
 PIN vss.gds716
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.542 8.1155 51.598 8.3155 ;
 END
 END vss.gds716
 PIN vss.gds717
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 7.9635 51.418 8.1635 ;
 END
 END vss.gds717
 PIN vss.gds718
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 7.8665 50.594 8.0665 ;
 END
 END vss.gds718
 PIN vss.gds719
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.09 7.843 52.13 8.043 ;
 END
 END vss.gds719
 PIN vss.gds720
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.47 8.0595 52.53 8.2595 ;
 END
 END vss.gds720
 PIN vss.gds721
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 7.981 52.362 8.181 ;
 END
 END vss.gds721
 PIN vss.gds722
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 50.624 9.176 50.68 9.329 ;
 RECT 50.624 6.656 50.68 6.809 ;
 RECT 50.624 7.916 50.68 8.069 ;
 RECT 50.624 10.436 50.68 10.589 ;
 RECT 50.456 7.5395 50.512 7.7395 ;
 RECT 50.96 7.2875 51.016 7.4875 ;
 RECT 50.456 8.7995 50.512 8.9995 ;
 RECT 50.96 8.5475 51.016 8.7475 ;
 RECT 50.96 6.0275 51.016 6.2275 ;
 RECT 50.456 6.2795 50.512 6.4795 ;
 RECT 50.456 10.0595 50.512 10.2595 ;
 RECT 50.96 9.8075 51.016 10.0075 ;
 RECT 51.968 7.954 52.024 8.154 ;
 RECT 51.8 7.9615 51.856 8.1615 ;
 RECT 51.632 7.954 51.688 8.154 ;
 RECT 51.464 7.954 51.52 8.154 ;
 RECT 51.296 7.954 51.352 8.154 ;
 RECT 52.136 7.954 52.192 8.154 ;
 RECT 51.128 8.069 51.184 8.269 ;
 END
 END vss.gds722
 PIN vss.gds723
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.946 8.0595 60.006 8.2595 ;
 END
 END vss.gds723
 PIN vss.gds724
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.778 8.0595 59.838 8.2595 ;
 END
 END vss.gds724
 PIN vss.gds725
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.61 8.0595 59.67 8.2595 ;
 END
 END vss.gds725
 PIN vss.gds726
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.274 8.0595 59.334 8.2595 ;
 END
 END vss.gds726
 PIN vss.gds727
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.106 8.0595 59.166 8.2595 ;
 END
 END vss.gds727
 PIN vss.gds728
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.938 8.0595 58.998 8.2595 ;
 END
 END vss.gds728
 PIN vss.gds729
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.602 8.0595 58.662 8.2595 ;
 END
 END vss.gds729
 PIN vss.gds730
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.434 8.0595 58.494 8.2595 ;
 END
 END vss.gds730
 PIN vss.gds731
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.266 8.0595 58.326 8.2595 ;
 END
 END vss.gds731
 PIN vss.gds732
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.326 8.0595 55.386 8.2595 ;
 END
 END vss.gds732
 PIN vss.gds733
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.494 8.0595 55.554 8.2595 ;
 END
 END vss.gds733
 PIN vss.gds734
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 8.0595 60.174 8.2595 ;
 END
 END vss.gds734
 PIN vss.gds735
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 8.0595 59.502 8.2595 ;
 END
 END vss.gds735
 PIN vss.gds736
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 8.0595 58.83 8.2595 ;
 END
 END vss.gds736
 PIN vss.gds737
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 8.0595 55.722 8.2595 ;
 END
 END vss.gds737
 PIN vss.gds738
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.83 8.0595 55.89 8.2595 ;
 END
 END vss.gds738
 PIN vss.gds739
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.998 8.0595 56.058 8.2595 ;
 END
 END vss.gds739
 PIN vss.gds740
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.166 8.0595 56.226 8.2595 ;
 END
 END vss.gds740
 PIN vss.gds741
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 8.0595 56.394 8.2595 ;
 END
 END vss.gds741
 PIN vss.gds742
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.502 8.0595 56.562 8.2595 ;
 END
 END vss.gds742
 PIN vss.gds743
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.67 8.0595 56.73 8.2595 ;
 END
 END vss.gds743
 PIN vss.gds744
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.838 8.0595 56.898 8.2595 ;
 END
 END vss.gds744
 PIN vss.gds745
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.342 8.0595 57.402 8.2595 ;
 END
 END vss.gds745
 PIN vss.gds746
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.51 8.0595 57.57 8.2595 ;
 END
 END vss.gds746
 PIN vss.gds747
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 8.0595 57.738 8.2595 ;
 END
 END vss.gds747
 PIN vss.gds748
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.174 8.0595 57.234 8.2595 ;
 END
 END vss.gds748
 PIN vss.gds749
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 8.0595 57.066 8.2595 ;
 END
 END vss.gds749
 PIN vss.gds750
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 58.016 9.896 58.072 10.096 ;
 RECT 58.016 7.376 58.072 7.576 ;
 RECT 58.016 8.636 58.072 8.836 ;
 RECT 58.016 6.116 58.072 6.316 ;
 RECT 57.848 8.006 57.904 8.206 ;
 END
 END vss.gds750
 PIN vss.gds751
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 8.978 65.054 9.178 ;
 END
 END vss.gds751
 PIN vss.gds752
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 6.458 65.054 6.658 ;
 END
 END vss.gds752
 PIN vss.gds753
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 7.718 65.054 7.918 ;
 END
 END vss.gds753
 PIN vss.gds754
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 10.238 65.054 10.438 ;
 END
 END vss.gds754
 PIN vss.gds755
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 8.1155 64.214 8.3155 ;
 END
 END vss.gds755
 PIN vss.gds756
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.418 8.112 64.474 8.312 ;
 END
 END vss.gds756
 PIN vss.gds757
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.306 8.0595 63.366 8.2595 ;
 END
 END vss.gds757
 PIN vss.gds758
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.138 8.0595 63.198 8.2595 ;
 END
 END vss.gds758
 PIN vss.gds759
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.97 8.0595 63.03 8.2595 ;
 END
 END vss.gds759
 PIN vss.gds760
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.634 8.0595 62.694 8.2595 ;
 END
 END vss.gds760
 PIN vss.gds761
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.466 8.0595 62.526 8.2595 ;
 END
 END vss.gds761
 PIN vss.gds762
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.298 8.0595 62.358 8.2595 ;
 END
 END vss.gds762
 PIN vss.gds763
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.962 8.0595 62.022 8.2595 ;
 END
 END vss.gds763
 PIN vss.gds764
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.794 8.0595 61.854 8.2595 ;
 END
 END vss.gds764
 PIN vss.gds765
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.626 8.0595 61.686 8.2595 ;
 END
 END vss.gds765
 PIN vss.gds766
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.29 8.0595 61.35 8.2595 ;
 END
 END vss.gds766
 PIN vss.gds767
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.122 8.0595 61.182 8.2595 ;
 END
 END vss.gds767
 PIN vss.gds768
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.954 8.0595 61.014 8.2595 ;
 END
 END vss.gds768
 PIN vss.gds769
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.618 8.0595 60.678 8.2595 ;
 END
 END vss.gds769
 PIN vss.gds770
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.45 8.0595 60.51 8.2595 ;
 END
 END vss.gds770
 PIN vss.gds771
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.282 8.0595 60.342 8.2595 ;
 END
 END vss.gds771
 PIN vss.gds772
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 7.981 63.534 8.181 ;
 END
 END vss.gds772
 PIN vss.gds773
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 8.0595 62.862 8.2595 ;
 END
 END vss.gds773
 PIN vss.gds774
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 8.0595 62.19 8.2595 ;
 END
 END vss.gds774
 PIN vss.gds775
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 8.0595 61.518 8.2595 ;
 END
 END vss.gds775
 PIN vss.gds776
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 8.0595 60.846 8.2595 ;
 END
 END vss.gds776
 PIN vss.gds777
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 7.9635 63.974 8.1635 ;
 END
 END vss.gds777
 PIN vss.gds778
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 7.843 63.746 8.043 ;
 END
 END vss.gds778
 PIN vss.gds779
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 8.0595 64.814 8.2595 ;
 END
 END vss.gds779
 PIN vss.gds780
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 65.156 9.156 65.212 9.329 ;
 RECT 65.156 6.636 65.212 6.809 ;
 RECT 65.156 7.896 65.212 8.069 ;
 RECT 65.156 10.416 65.212 10.589 ;
 RECT 64.82 9.883 64.876 10.083 ;
 RECT 64.82 7.363 64.876 7.563 ;
 RECT 64.82 6.103 64.876 6.303 ;
 RECT 64.82 8.623 64.876 8.823 ;
 RECT 64.652 7.935 64.708 8.135 ;
 RECT 64.484 7.873 64.54 8.073 ;
 RECT 64.316 7.924 64.372 8.124 ;
 RECT 64.148 7.924 64.204 8.124 ;
 RECT 63.98 7.924 64.036 8.124 ;
 RECT 63.644 7.954 63.7 8.154 ;
 RECT 63.812 7.954 63.868 8.154 ;
 END
 END vss.gds780
 PIN vss.gds781
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 7.758 66.026 7.958 ;
 END
 END vss.gds781
 PIN vss.gds782
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 6.498 66.026 6.698 ;
 END
 END vss.gds782
 PIN vss.gds783
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 9.018 66.026 9.218 ;
 END
 END vss.gds783
 PIN vss.gds784
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 10.278 66.026 10.478 ;
 END
 END vss.gds784
 PIN vss.gds785
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.69 8.0595 69.75 8.2595 ;
 END
 END vss.gds785
 PIN vss.gds786
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.858 8.0595 69.918 8.2595 ;
 END
 END vss.gds786
 PIN vss.gds787
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.194 8.0595 70.254 8.2595 ;
 END
 END vss.gds787
 PIN vss.gds788
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 8.0185 68.15 8.2185 ;
 END
 END vss.gds788
 PIN vss.gds789
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 8.1 66.318 8.3 ;
 END
 END vss.gds789
 PIN vss.gds790
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 8.0595 70.086 8.2595 ;
 END
 END vss.gds790
 PIN vss.gds791
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 8.1 66.998 8.3 ;
 END
 END vss.gds791
 PIN vss.gds792
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 8.1 65.654 8.3 ;
 END
 END vss.gds792
 PIN vss.gds793
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 7.8665 67.646 8.0665 ;
 END
 END vss.gds793
 PIN vss.gds794
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 7.956 66.574 8.156 ;
 END
 END vss.gds794
 PIN vss.gds795
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 8.112 67.97 8.312 ;
 END
 END vss.gds795
 PIN vss.gds796
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 8.473 67.302 8.673 ;
 END
 END vss.gds796
 PIN vss.gds797
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 9.733 67.302 9.933 ;
 END
 END vss.gds797
 PIN vss.gds798
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 7.213 67.302 7.413 ;
 END
 END vss.gds798
 PIN vss.gds799
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 5.953 67.302 6.153 ;
 END
 END vss.gds799
 PIN vss.gds800
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 7.9635 68.99 8.1635 ;
 END
 END vss.gds800
 PIN vss.gds801
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.594 8.1155 68.65 8.3155 ;
 END
 END vss.gds801
 PIN vss.gds802
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 7.9635 68.47 8.1635 ;
 END
 END vss.gds802
 PIN vss.gds803
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.142 7.843 69.182 8.043 ;
 END
 END vss.gds803
 PIN vss.gds804
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.522 8.0595 69.582 8.2595 ;
 END
 END vss.gds804
 PIN vss.gds805
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 7.981 69.414 8.181 ;
 END
 END vss.gds805
 PIN vss.gds806
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 67.676 9.176 67.732 9.329 ;
 RECT 65.324 9.129 65.38 9.329 ;
 RECT 66.92 9.173 66.976 9.338 ;
 RECT 66.752 9.173 66.808 9.338 ;
 RECT 65.996 9.173 66.052 9.338 ;
 RECT 65.828 9.173 65.884 9.338 ;
 RECT 67.676 6.656 67.732 6.809 ;
 RECT 65.324 6.609 65.38 6.809 ;
 RECT 66.92 6.653 66.976 6.818 ;
 RECT 66.752 6.653 66.808 6.818 ;
 RECT 65.996 6.653 66.052 6.818 ;
 RECT 65.828 6.653 65.884 6.818 ;
 RECT 66.752 9.4 66.808 9.6 ;
 RECT 67.004 9.403 67.06 9.603 ;
 RECT 67.676 7.916 67.732 8.069 ;
 RECT 65.324 7.869 65.38 8.069 ;
 RECT 66.92 7.913 66.976 8.078 ;
 RECT 66.752 7.913 66.808 8.078 ;
 RECT 65.996 7.913 66.052 8.078 ;
 RECT 65.828 7.913 65.884 8.078 ;
 RECT 67.676 10.436 67.732 10.589 ;
 RECT 65.324 10.389 65.38 10.589 ;
 RECT 66.92 10.433 66.976 10.598 ;
 RECT 66.752 10.433 66.808 10.598 ;
 RECT 65.996 10.433 66.052 10.598 ;
 RECT 65.828 10.433 65.884 10.598 ;
 RECT 66.752 5.62 66.808 5.82 ;
 RECT 67.004 5.623 67.06 5.823 ;
 RECT 66.752 6.88 66.808 7.08 ;
 RECT 67.004 6.883 67.06 7.083 ;
 RECT 66.752 8.14 66.808 8.34 ;
 RECT 67.004 8.143 67.06 8.343 ;
 RECT 66.164 9.959 66.22 10.159 ;
 RECT 65.492 9.749 65.548 9.949 ;
 RECT 65.324 9.749 65.38 9.949 ;
 RECT 67.508 10.0595 67.564 10.2595 ;
 RECT 68.012 9.8075 68.068 10.0075 ;
 RECT 66.584 9.959 66.64 10.159 ;
 RECT 65.492 8.489 65.548 8.689 ;
 RECT 65.324 8.489 65.38 8.689 ;
 RECT 67.508 8.7995 67.564 8.9995 ;
 RECT 68.012 8.5475 68.068 8.7475 ;
 RECT 66.164 7.439 66.22 7.639 ;
 RECT 65.492 7.229 65.548 7.429 ;
 RECT 65.324 7.229 65.38 7.429 ;
 RECT 67.508 7.5395 67.564 7.7395 ;
 RECT 68.012 7.2875 68.068 7.4875 ;
 RECT 66.584 7.439 66.64 7.639 ;
 RECT 68.012 6.0275 68.068 6.2275 ;
 RECT 67.508 6.2795 67.564 6.4795 ;
 RECT 66.164 6.179 66.22 6.379 ;
 RECT 66.584 6.179 66.64 6.379 ;
 RECT 65.492 5.969 65.548 6.169 ;
 RECT 65.324 5.969 65.38 6.169 ;
 RECT 66.164 8.699 66.22 8.899 ;
 RECT 66.584 8.699 66.64 8.899 ;
 RECT 66.332 8.1395 66.388 8.3395 ;
 RECT 69.02 7.954 69.076 8.154 ;
 RECT 68.852 7.9615 68.908 8.1615 ;
 RECT 68.684 7.954 68.74 8.154 ;
 RECT 68.516 7.954 68.572 8.154 ;
 RECT 68.348 7.954 68.404 8.154 ;
 RECT 69.188 7.954 69.244 8.154 ;
 RECT 68.18 8.069 68.236 8.269 ;
 END
 END vss.gds806
 PIN vss.gds807
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.362 8.0595 70.422 8.2595 ;
 END
 END vss.gds807
 PIN vss.gds808
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.53 8.0595 70.59 8.2595 ;
 END
 END vss.gds808
 PIN vss.gds809
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.866 8.0595 70.926 8.2595 ;
 END
 END vss.gds809
 PIN vss.gds810
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.034 8.0595 71.094 8.2595 ;
 END
 END vss.gds810
 PIN vss.gds811
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.202 8.0595 71.262 8.2595 ;
 END
 END vss.gds811
 PIN vss.gds812
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.538 8.0595 71.598 8.2595 ;
 END
 END vss.gds812
 PIN vss.gds813
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.706 8.0595 71.766 8.2595 ;
 END
 END vss.gds813
 PIN vss.gds814
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.874 8.0595 71.934 8.2595 ;
 END
 END vss.gds814
 PIN vss.gds815
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.21 8.0595 72.27 8.2595 ;
 END
 END vss.gds815
 PIN vss.gds816
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.378 8.0595 72.438 8.2595 ;
 END
 END vss.gds816
 PIN vss.gds817
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.546 8.0595 72.606 8.2595 ;
 END
 END vss.gds817
 PIN vss.gds818
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.882 8.0595 72.942 8.2595 ;
 END
 END vss.gds818
 PIN vss.gds819
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.05 8.0595 73.11 8.2595 ;
 END
 END vss.gds819
 PIN vss.gds820
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 8.0595 71.43 8.2595 ;
 END
 END vss.gds820
 PIN vss.gds821
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 8.0595 72.102 8.2595 ;
 END
 END vss.gds821
 PIN vss.gds822
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 8.0595 72.774 8.2595 ;
 END
 END vss.gds822
 PIN vss.gds823
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 8.0595 70.758 8.2595 ;
 END
 END vss.gds823
 PIN vss.gds824
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.554 8.0595 73.614 8.2595 ;
 END
 END vss.gds824
 PIN vss.gds825
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.722 8.0595 73.782 8.2595 ;
 END
 END vss.gds825
 PIN vss.gds826
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 8.0595 73.446 8.2595 ;
 END
 END vss.gds826
 PIN vss.gds827
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.218 8.0595 73.278 8.2595 ;
 END
 END vss.gds827
 PIN vss.gds828
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.89 8.0595 73.95 8.2595 ;
 END
 END vss.gds828
 PIN vss.gds829
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.394 8.0595 74.454 8.2595 ;
 END
 END vss.gds829
 PIN vss.gds830
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 8.0595 74.118 8.2595 ;
 END
 END vss.gds830
 PIN vss.gds831
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.562 8.0595 74.622 8.2595 ;
 END
 END vss.gds831
 PIN vss.gds832
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 8.0595 74.79 8.2595 ;
 END
 END vss.gds832
 PIN vss.gds833
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.226 8.0595 74.286 8.2595 ;
 END
 END vss.gds833
 PIN vss.gds834
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 10.993 2.962 11.193 ;
 END
 END vss.gds834
 PIN vss.gds835
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 12.253 2.962 12.453 ;
 END
 END vss.gds835
 PIN vss.gds836
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 13.513 2.962 13.713 ;
 END
 END vss.gds836
 PIN vss.gds837
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 14.773 2.962 14.973 ;
 END
 END vss.gds837
 PIN vss.gds838
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 11.852 3.142 12.052 ;
 END
 END vss.gds838
 PIN vss.gds839
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 10.592 3.142 10.792 ;
 END
 END vss.gds839
 PIN vss.gds840
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 14.372 3.142 14.572 ;
 END
 END vss.gds840
 PIN vss.gds841
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 12.477 0.942 12.677 ;
 END
 END vss.gds841
 PIN vss.gds842
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.286 12.883 3.326 13.083 ;
 END
 END vss.gds842
 PIN vss.gds843
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 12.883 4.194 13.083 ;
 END
 END vss.gds843
 PIN vss.gds844
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 13.112 3.142 13.312 ;
 END
 END vss.gds844
 PIN vss.gds845
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 12.883 5.074 13.083 ;
 END
 END vss.gds845
 PIN vss.gds846
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 12.5775 0.718 12.7775 ;
 END
 END vss.gds846
 PIN vss.gds847
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.442 12.477 4.482 12.677 ;
 END
 END vss.gds847
 PIN vss.gds848
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.57 12.68 4.61 12.88 ;
 END
 END vss.gds848
 PIN vss.gds849
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 12.477 4.882 12.677 ;
 END
 END vss.gds849
 PIN vss.gds850
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 12.678 0.602 12.878 ;
 END
 END vss.gds850
 PIN vss.gds851
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 12.9065 2.122 13.1065 ;
 END
 END vss.gds851
 PIN vss.gds852
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 13.021 1.282 13.221 ;
 END
 END vss.gds852
 PIN vss.gds853
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 13.2555 1.462 13.4555 ;
 END
 END vss.gds853
 PIN vss.gds854
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.414 13.159 3.454 13.359 ;
 END
 END vss.gds854
 PIN vss.gds855
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.562 13.159 3.602 13.359 ;
 END
 END vss.gds855
 PIN vss.gds856
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 12.818 2.302 13.018 ;
 END
 END vss.gds856
 PIN vss.gds857
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 12.7795 4.002 12.9795 ;
 END
 END vss.gds857
 PIN vss.gds858
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 12.7795 5.282 12.9795 ;
 END
 END vss.gds858
 PIN vss.gds859
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 12.8115 0.29 13.0115 ;
 END
 END vss.gds859
 PIN vss.gds860
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.754 12.883 3.794 13.083 ;
 END
 END vss.gds860
 PIN vss.gds861
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 2.576 10.9935 2.632 11.1935 ;
 RECT 2.408 10.9935 2.464 11.1935 ;
 RECT 2.996 10.9935 3.052 11.1935 ;
 RECT 3.332 11.085 3.388 11.285 ;
 RECT 2.408 12.2535 2.464 12.4535 ;
 RECT 2.576 12.2535 2.632 12.4535 ;
 RECT 2.996 12.2535 3.052 12.4535 ;
 RECT 3.332 12.345 3.388 12.545 ;
 RECT 3.5 12.3015 3.556 12.5015 ;
 RECT 0.98 12.1685 1.036 12.3685 ;
 RECT 2.072 12.169 2.128 12.369 ;
 RECT 0.812 11.085 0.868 11.285 ;
 RECT 3.752 13.789 3.808 13.989 ;
 RECT 3.5 13.5615 3.556 13.7615 ;
 RECT 0.98 13.4285 1.036 13.6285 ;
 RECT 2.576 13.5135 2.632 13.7135 ;
 RECT 2.072 13.429 2.128 13.629 ;
 RECT 2.408 13.5135 2.464 13.7135 ;
 RECT 2.996 13.5135 3.052 13.7135 ;
 RECT 2.744 13.429 2.8 13.629 ;
 RECT 3.332 13.605 3.388 13.805 ;
 RECT 3.164 13.519 3.22 13.719 ;
 RECT 2.408 14.7735 2.464 14.9735 ;
 RECT 2.576 14.7735 2.632 14.9735 ;
 RECT 2.996 14.7735 3.052 14.9735 ;
 RECT 3.332 14.865 3.388 15.065 ;
 RECT 3.5 14.8215 3.556 15.0215 ;
 RECT 0.98 14.6885 1.036 14.8885 ;
 RECT 2.072 14.689 2.128 14.889 ;
 RECT 0.392 13.519 0.448 13.719 ;
 RECT 0.812 13.605 0.868 13.805 ;
 RECT 0.644 13.519 0.7 13.719 ;
 RECT 1.232 13.519 1.288 13.719 ;
 RECT 1.4 13.519 1.456 13.719 ;
 RECT 1.568 13.519 1.624 13.719 ;
 RECT 1.82 13.519 1.876 13.719 ;
 RECT 2.24 13.519 2.296 13.719 ;
 RECT 0.392 14.779 0.448 14.979 ;
 RECT 0.812 14.865 0.868 15.065 ;
 RECT 0.644 14.779 0.7 14.979 ;
 RECT 1.232 14.779 1.288 14.979 ;
 RECT 1.4 14.779 1.456 14.979 ;
 RECT 1.568 14.779 1.624 14.979 ;
 RECT 1.82 14.779 1.876 14.979 ;
 RECT 2.24 14.779 2.296 14.979 ;
 RECT 2.744 14.689 2.8 14.889 ;
 RECT 3.164 14.779 3.22 14.979 ;
 RECT 3.92 14.779 3.976 14.979 ;
 RECT 3.752 15.049 3.808 15.249 ;
 RECT 4.508 14.9785 4.564 15.1785 ;
 RECT 4.508 13.7185 4.564 13.9185 ;
 RECT 3.92 13.519 3.976 13.719 ;
 RECT 3.5 11.0415 3.556 11.2415 ;
 RECT 0.392 10.999 0.448 11.199 ;
 RECT 0.644 10.999 0.7 11.199 ;
 RECT 1.232 10.999 1.288 11.199 ;
 RECT 0.98 10.9085 1.036 11.1085 ;
 RECT 1.4 10.999 1.456 11.199 ;
 RECT 1.568 10.999 1.624 11.199 ;
 RECT 2.072 10.909 2.128 11.109 ;
 RECT 1.82 10.999 1.876 11.199 ;
 RECT 2.744 10.909 2.8 11.109 ;
 RECT 3.164 10.999 3.22 11.199 ;
 RECT 2.24 10.999 2.296 11.199 ;
 RECT 0.392 12.259 0.448 12.459 ;
 RECT 0.812 12.345 0.868 12.545 ;
 RECT 0.644 12.259 0.7 12.459 ;
 RECT 1.232 12.259 1.288 12.459 ;
 RECT 1.4 12.259 1.456 12.459 ;
 RECT 1.568 12.259 1.624 12.459 ;
 RECT 1.82 12.259 1.876 12.459 ;
 RECT 2.24 12.259 2.296 12.459 ;
 RECT 2.744 12.169 2.8 12.369 ;
 RECT 3.164 12.259 3.22 12.459 ;
 RECT 3.92 12.259 3.976 12.459 ;
 RECT 3.752 12.529 3.808 12.729 ;
 RECT 4.508 12.4585 4.564 12.6585 ;
 RECT 3.92 10.999 3.976 11.199 ;
 RECT 3.752 11.269 3.808 11.469 ;
 RECT 4.508 11.1985 4.564 11.3985 ;
 END
 END vss.gds861
 PIN vss.gds862
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.134 13.0995 10.194 13.2995 ;
 END
 END vss.gds862
 PIN vss.gds863
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.966 13.0995 10.026 13.2995 ;
 END
 END vss.gds863
 PIN vss.gds864
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.798 13.0995 9.858 13.2995 ;
 END
 END vss.gds864
 PIN vss.gds865
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 13.0995 9.69 13.2995 ;
 END
 END vss.gds865
 PIN vss.gds866
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.462 13.0995 9.522 13.2995 ;
 END
 END vss.gds866
 PIN vss.gds867
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 13.0995 9.018 13.2995 ;
 END
 END vss.gds867
 PIN vss.gds868
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.79 13.0995 8.85 13.2995 ;
 END
 END vss.gds868
 PIN vss.gds869
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.622 13.0995 8.682 13.2995 ;
 END
 END vss.gds869
 PIN vss.gds870
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.454 13.0995 8.514 13.2995 ;
 END
 END vss.gds870
 PIN vss.gds871
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 12.883 5.474 13.083 ;
 END
 END vss.gds871
 PIN vss.gds872
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 13.0995 8.346 13.2995 ;
 END
 END vss.gds872
 PIN vss.gds873
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.118 13.0995 8.178 13.2995 ;
 END
 END vss.gds873
 PIN vss.gds874
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.95 13.0995 8.01 13.2995 ;
 END
 END vss.gds874
 PIN vss.gds875
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.294 13.0995 9.354 13.2995 ;
 END
 END vss.gds875
 PIN vss.gds876
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.782 13.0995 7.842 13.2995 ;
 END
 END vss.gds876
 PIN vss.gds877
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 13.0995 7.674 13.2995 ;
 END
 END vss.gds877
 PIN vss.gds878
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.126 13.0995 9.186 13.2995 ;
 END
 END vss.gds878
 PIN vss.gds879
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.446 13.0995 7.506 13.2995 ;
 END
 END vss.gds879
 PIN vss.gds880
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.278 13.0995 7.338 13.2995 ;
 END
 END vss.gds880
 PIN vss.gds881
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.11 13.0995 7.17 13.2995 ;
 END
 END vss.gds881
 PIN vss.gds882
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 12.883 5.73 13.083 ;
 END
 END vss.gds882
 PIN vss.gds883
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 12.883 5.986 13.083 ;
 END
 END vss.gds883
 PIN vss.gds884
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 12.679 6.434 12.879 ;
 END
 END vss.gds884
 PIN vss.gds885
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 12.68 6.178 12.88 ;
 END
 END vss.gds885
 PIN vss.gds886
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 6.608 15.049 6.664 15.249 ;
 RECT 6.524 14.772 6.58 14.972 ;
 RECT 6.692 14.922 6.748 15.122 ;
 RECT 6.692 13.662 6.748 13.862 ;
 RECT 6.524 13.512 6.58 13.712 ;
 RECT 6.608 13.789 6.664 13.989 ;
 RECT 6.608 12.529 6.664 12.729 ;
 RECT 6.524 12.252 6.58 12.452 ;
 RECT 6.692 12.402 6.748 12.602 ;
 RECT 6.692 11.142 6.748 11.342 ;
 RECT 6.524 10.992 6.58 11.192 ;
 RECT 6.608 11.269 6.664 11.469 ;
 END
 END vss.gds886
 PIN vss.gds887
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 12.758 13.898 12.958 ;
 END
 END vss.gds887
 PIN vss.gds888
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 12.798 14.87 12.998 ;
 END
 END vss.gds888
 PIN vss.gds889
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 11.498 13.898 11.698 ;
 END
 END vss.gds889
 PIN vss.gds890
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 11.538 14.87 11.738 ;
 END
 END vss.gds890
 PIN vss.gds891
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 14.018 13.898 14.218 ;
 END
 END vss.gds891
 PIN vss.gds892
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 14.058 14.87 14.258 ;
 END
 END vss.gds892
 PIN vss.gds893
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 15.278 13.898 15.478 ;
 END
 END vss.gds893
 PIN vss.gds894
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 15.318 14.87 15.518 ;
 END
 END vss.gds894
 PIN vss.gds895
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.15 13.0995 12.21 13.2995 ;
 END
 END vss.gds895
 PIN vss.gds896
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.982 13.0995 12.042 13.2995 ;
 END
 END vss.gds896
 PIN vss.gds897
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.814 13.0995 11.874 13.2995 ;
 END
 END vss.gds897
 PIN vss.gds898
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.478 13.0995 11.538 13.2995 ;
 END
 END vss.gds898
 PIN vss.gds899
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.31 13.0995 11.37 13.2995 ;
 END
 END vss.gds899
 PIN vss.gds900
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 13.1555 13.058 13.3555 ;
 END
 END vss.gds900
 PIN vss.gds901
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 13.0995 11.706 13.2995 ;
 END
 END vss.gds901
 PIN vss.gds902
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.142 13.0995 11.202 13.2995 ;
 END
 END vss.gds902
 PIN vss.gds903
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.806 13.0995 10.866 13.2995 ;
 END
 END vss.gds903
 PIN vss.gds904
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.638 13.0995 10.698 13.2995 ;
 END
 END vss.gds904
 PIN vss.gds905
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.47 13.0995 10.53 13.2995 ;
 END
 END vss.gds905
 PIN vss.gds906
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 13.0995 11.034 13.2995 ;
 END
 END vss.gds906
 PIN vss.gds907
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 13.0995 10.362 13.2995 ;
 END
 END vss.gds907
 PIN vss.gds908
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 13.14 15.162 13.34 ;
 END
 END vss.gds908
 PIN vss.gds909
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 13.14 14.498 13.34 ;
 END
 END vss.gds909
 PIN vss.gds910
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 13.0995 13.658 13.2995 ;
 END
 END vss.gds910
 PIN vss.gds911
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.262 13.152 13.318 13.352 ;
 END
 END vss.gds911
 PIN vss.gds912
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 13.021 12.378 13.221 ;
 END
 END vss.gds912
 PIN vss.gds913
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 12.883 12.59 13.083 ;
 END
 END vss.gds913
 PIN vss.gds914
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 13.0035 12.818 13.2035 ;
 END
 END vss.gds914
 PIN vss.gds915
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 14 14.196 14.056 14.369 ;
 RECT 14.168 14.169 14.224 14.369 ;
 RECT 14 11.676 14.056 11.849 ;
 RECT 14.168 11.649 14.224 11.849 ;
 RECT 14 12.936 14.056 13.109 ;
 RECT 14.168 12.909 14.224 13.109 ;
 RECT 14 15.456 14.056 15.629 ;
 RECT 14.168 15.429 14.224 15.629 ;
 RECT 14.336 12.269 14.392 12.469 ;
 RECT 14.168 12.269 14.224 12.469 ;
 RECT 14.336 11.009 14.392 11.209 ;
 RECT 14.168 11.009 14.224 11.209 ;
 RECT 14.336 13.529 14.392 13.729 ;
 RECT 14.168 13.529 14.224 13.729 ;
 RECT 14.336 14.789 14.392 14.989 ;
 RECT 14.168 14.789 14.224 14.989 ;
 RECT 13.664 14.923 13.72 15.123 ;
 RECT 15.008 14.999 15.064 15.199 ;
 RECT 14.84 15.473 14.896 15.638 ;
 RECT 14.672 15.473 14.728 15.638 ;
 RECT 13.664 12.403 13.72 12.603 ;
 RECT 15.008 12.479 15.064 12.679 ;
 RECT 14.84 12.953 14.896 13.118 ;
 RECT 14.672 12.953 14.728 13.118 ;
 RECT 13.664 11.143 13.72 11.343 ;
 RECT 15.008 11.219 15.064 11.419 ;
 RECT 14.84 11.693 14.896 11.858 ;
 RECT 14.672 11.693 14.728 11.858 ;
 RECT 15.008 13.739 15.064 13.939 ;
 RECT 14.84 14.213 14.896 14.378 ;
 RECT 14.672 14.213 14.728 14.378 ;
 RECT 13.664 13.663 13.72 13.863 ;
 RECT 15.176 13.1795 15.232 13.3795 ;
 RECT 12.824 12.964 12.88 13.164 ;
 RECT 13.496 12.975 13.552 13.175 ;
 RECT 12.488 12.994 12.544 13.194 ;
 RECT 13.328 12.913 13.384 13.113 ;
 RECT 13.16 12.964 13.216 13.164 ;
 RECT 12.992 12.964 13.048 13.164 ;
 RECT 12.656 12.994 12.712 13.194 ;
 END
 END vss.gds915
 PIN vss.gds916
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 10.993 16.146 11.193 ;
 END
 END vss.gds916
 PIN vss.gds917
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 13.513 16.146 13.713 ;
 END
 END vss.gds917
 PIN vss.gds918
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 12.996 15.418 13.196 ;
 END
 END vss.gds918
 PIN vss.gds919
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 13.0995 20.274 13.2995 ;
 END
 END vss.gds919
 PIN vss.gds920
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 13.0995 18.93 13.2995 ;
 END
 END vss.gds920
 PIN vss.gds921
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.038 13.0995 19.098 13.2995 ;
 END
 END vss.gds921
 PIN vss.gds922
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.206 13.0995 19.266 13.2995 ;
 END
 END vss.gds922
 PIN vss.gds923
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.374 13.0995 19.434 13.2995 ;
 END
 END vss.gds923
 PIN vss.gds924
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 13.0995 19.602 13.2995 ;
 END
 END vss.gds924
 PIN vss.gds925
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 13.0035 17.314 13.2035 ;
 END
 END vss.gds925
 PIN vss.gds926
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 13.0585 16.994 13.2585 ;
 END
 END vss.gds926
 PIN vss.gds927
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 14.773 16.146 14.973 ;
 END
 END vss.gds927
 PIN vss.gds928
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.71 13.0995 19.77 13.2995 ;
 END
 END vss.gds928
 PIN vss.gds929
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.878 13.0995 19.938 13.2995 ;
 END
 END vss.gds929
 PIN vss.gds930
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 12.253 16.146 12.453 ;
 END
 END vss.gds930
 PIN vss.gds931
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 13.14 15.842 13.34 ;
 END
 END vss.gds931
 PIN vss.gds932
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 13.152 16.814 13.352 ;
 END
 END vss.gds932
 PIN vss.gds933
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.046 13.0995 20.106 13.2995 ;
 END
 END vss.gds933
 PIN vss.gds934
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.702 13.0995 18.762 13.2995 ;
 END
 END vss.gds934
 PIN vss.gds935
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.534 13.0995 18.594 13.2995 ;
 END
 END vss.gds935
 PIN vss.gds936
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.366 13.0995 18.426 13.2995 ;
 END
 END vss.gds936
 PIN vss.gds937
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 13.021 18.258 13.221 ;
 END
 END vss.gds937
 PIN vss.gds938
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 13.0035 17.834 13.2035 ;
 END
 END vss.gds938
 PIN vss.gds939
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.438 13.1555 17.494 13.3555 ;
 END
 END vss.gds939
 PIN vss.gds940
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 12.9065 16.49 13.1065 ;
 END
 END vss.gds940
 PIN vss.gds941
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.986 12.883 18.026 13.083 ;
 END
 END vss.gds941
 PIN vss.gds942
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 15.596 13.18 15.652 13.38 ;
 RECT 15.848 13.183 15.904 13.383 ;
 RECT 16.52 14.216 16.576 14.369 ;
 RECT 15.764 14.213 15.82 14.378 ;
 RECT 15.596 14.213 15.652 14.378 ;
 RECT 15.596 10.66 15.652 10.86 ;
 RECT 15.848 10.663 15.904 10.863 ;
 RECT 16.52 11.696 16.576 11.849 ;
 RECT 15.764 11.693 15.82 11.858 ;
 RECT 15.596 11.693 15.652 11.858 ;
 RECT 15.596 11.92 15.652 12.12 ;
 RECT 15.848 11.923 15.904 12.123 ;
 RECT 16.52 12.956 16.576 13.109 ;
 RECT 15.764 12.953 15.82 13.118 ;
 RECT 15.596 12.953 15.652 13.118 ;
 RECT 15.596 14.44 15.652 14.64 ;
 RECT 15.848 14.443 15.904 14.643 ;
 RECT 16.52 15.476 16.576 15.629 ;
 RECT 15.764 15.473 15.82 15.638 ;
 RECT 15.596 15.473 15.652 15.638 ;
 RECT 16.352 15.0995 16.408 15.2995 ;
 RECT 16.856 14.8475 16.912 15.0475 ;
 RECT 16.856 12.3275 16.912 12.5275 ;
 RECT 16.352 12.5795 16.408 12.7795 ;
 RECT 16.352 11.3195 16.408 11.5195 ;
 RECT 16.856 11.0675 16.912 11.2675 ;
 RECT 15.428 14.999 15.484 15.199 ;
 RECT 15.428 12.479 15.484 12.679 ;
 RECT 15.428 11.219 15.484 11.419 ;
 RECT 15.428 13.739 15.484 13.939 ;
 RECT 16.352 13.8395 16.408 14.0395 ;
 RECT 16.856 13.5875 16.912 13.7875 ;
 RECT 17.864 12.994 17.92 13.194 ;
 RECT 17.696 13.0015 17.752 13.2015 ;
 RECT 17.528 12.994 17.584 13.194 ;
 RECT 17.36 12.994 17.416 13.194 ;
 RECT 17.192 12.994 17.248 13.194 ;
 RECT 18.032 12.994 18.088 13.194 ;
 RECT 17.024 13.109 17.08 13.309 ;
 END
 END vss.gds942
 PIN vss.gds943
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.17 13.0995 25.23 13.2995 ;
 END
 END vss.gds943
 PIN vss.gds944
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.002 13.0995 25.062 13.2995 ;
 END
 END vss.gds944
 PIN vss.gds945
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.834 13.0995 24.894 13.2995 ;
 END
 END vss.gds945
 PIN vss.gds946
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.498 13.0995 24.558 13.2995 ;
 END
 END vss.gds946
 PIN vss.gds947
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.33 13.0995 24.39 13.2995 ;
 END
 END vss.gds947
 PIN vss.gds948
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.162 13.0995 24.222 13.2995 ;
 END
 END vss.gds948
 PIN vss.gds949
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.382 13.0995 20.442 13.2995 ;
 END
 END vss.gds949
 PIN vss.gds950
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.55 13.0995 20.61 13.2995 ;
 END
 END vss.gds950
 PIN vss.gds951
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.718 13.0995 20.778 13.2995 ;
 END
 END vss.gds951
 PIN vss.gds952
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.054 13.0995 21.114 13.2995 ;
 END
 END vss.gds952
 PIN vss.gds953
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.222 13.0995 21.282 13.2995 ;
 END
 END vss.gds953
 PIN vss.gds954
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.39 13.0995 21.45 13.2995 ;
 END
 END vss.gds954
 PIN vss.gds955
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.726 13.0995 21.786 13.2995 ;
 END
 END vss.gds955
 PIN vss.gds956
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.894 13.0995 21.954 13.2995 ;
 END
 END vss.gds956
 PIN vss.gds957
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.062 13.0995 22.122 13.2995 ;
 END
 END vss.gds957
 PIN vss.gds958
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.398 13.0995 22.458 13.2995 ;
 END
 END vss.gds958
 PIN vss.gds959
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.566 13.0995 22.626 13.2995 ;
 END
 END vss.gds959
 PIN vss.gds960
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.734 13.0995 22.794 13.2995 ;
 END
 END vss.gds960
 PIN vss.gds961
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 13.0995 24.726 13.2995 ;
 END
 END vss.gds961
 PIN vss.gds962
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 13.0995 21.618 13.2995 ;
 END
 END vss.gds962
 PIN vss.gds963
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 13.0995 20.946 13.2995 ;
 END
 END vss.gds963
 PIN vss.gds964
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 13.0995 22.29 13.2995 ;
 END
 END vss.gds964
 PIN vss.gds965
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 13.0995 22.962 13.2995 ;
 END
 END vss.gds965
 PIN vss.gds966
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.07 13.0995 23.13 13.2995 ;
 END
 END vss.gds966
 PIN vss.gds967
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.238 13.0995 23.298 13.2995 ;
 END
 END vss.gds967
 PIN vss.gds968
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.406 13.0995 23.466 13.2995 ;
 END
 END vss.gds968
 PIN vss.gds969
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 13.0995 23.634 13.2995 ;
 END
 END vss.gds969
 PIN vss.gds970
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 23.912 14.936 23.968 15.136 ;
 RECT 23.912 12.416 23.968 12.616 ;
 RECT 23.912 11.156 23.968 11.356 ;
 RECT 23.912 13.676 23.968 13.876 ;
 RECT 23.744 13.046 23.8 13.246 ;
 END
 END vss.gds970
 PIN vss.gds971
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.202 13.0995 29.262 13.2995 ;
 END
 END vss.gds971
 PIN vss.gds972
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.034 13.0995 29.094 13.2995 ;
 END
 END vss.gds972
 PIN vss.gds973
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.866 13.0995 28.926 13.2995 ;
 END
 END vss.gds973
 PIN vss.gds974
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.53 13.0995 28.59 13.2995 ;
 END
 END vss.gds974
 PIN vss.gds975
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.362 13.0995 28.422 13.2995 ;
 END
 END vss.gds975
 PIN vss.gds976
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.194 13.0995 28.254 13.2995 ;
 END
 END vss.gds976
 PIN vss.gds977
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.858 13.0995 27.918 13.2995 ;
 END
 END vss.gds977
 PIN vss.gds978
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.69 13.0995 27.75 13.2995 ;
 END
 END vss.gds978
 PIN vss.gds979
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.522 13.0995 27.582 13.2995 ;
 END
 END vss.gds979
 PIN vss.gds980
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.186 13.0995 27.246 13.2995 ;
 END
 END vss.gds980
 PIN vss.gds981
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.018 13.0995 27.078 13.2995 ;
 END
 END vss.gds981
 PIN vss.gds982
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.85 13.0995 26.91 13.2995 ;
 END
 END vss.gds982
 PIN vss.gds983
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.514 13.0995 26.574 13.2995 ;
 END
 END vss.gds983
 PIN vss.gds984
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.346 13.0995 26.406 13.2995 ;
 END
 END vss.gds984
 PIN vss.gds985
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.178 13.0995 26.238 13.2995 ;
 END
 END vss.gds985
 PIN vss.gds986
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.842 13.0995 25.902 13.2995 ;
 END
 END vss.gds986
 PIN vss.gds987
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.674 13.0995 25.734 13.2995 ;
 END
 END vss.gds987
 PIN vss.gds988
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.506 13.0995 25.566 13.2995 ;
 END
 END vss.gds988
 PIN vss.gds989
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 13.0995 28.758 13.2995 ;
 END
 END vss.gds989
 PIN vss.gds990
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 13.0995 28.086 13.2995 ;
 END
 END vss.gds990
 PIN vss.gds991
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 13.0995 27.414 13.2995 ;
 END
 END vss.gds991
 PIN vss.gds992
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 13.0995 26.742 13.2995 ;
 END
 END vss.gds992
 PIN vss.gds993
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 13.0995 26.07 13.2995 ;
 END
 END vss.gds993
 PIN vss.gds994
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 13.0995 25.398 13.2995 ;
 END
 END vss.gds994
 PIN vss.gds995
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 13.021 29.43 13.221 ;
 END
 END vss.gds995
 PIN vss.gds996
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 13.1555 30.11 13.3555 ;
 END
 END vss.gds996
 PIN vss.gds997
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 13.0035 29.87 13.2035 ;
 END
 END vss.gds997
 PIN vss.gds998
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 12.883 29.642 13.083 ;
 END
 END vss.gds998
 PIN vss.gds999
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.876 12.964 29.932 13.164 ;
 RECT 30.212 12.964 30.268 13.164 ;
 RECT 29.54 12.994 29.596 13.194 ;
 RECT 30.044 12.964 30.1 13.164 ;
 RECT 29.708 12.994 29.764 13.194 ;
 END
 END vss.gds999
 PIN vss.gds1000
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 12.798 31.922 12.998 ;
 END
 END vss.gds1000
 PIN vss.gds1001
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 11.498 30.95 11.698 ;
 END
 END vss.gds1001
 PIN vss.gds1002
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 11.538 31.922 11.738 ;
 END
 END vss.gds1002
 PIN vss.gds1003
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 14.058 31.922 14.258 ;
 END
 END vss.gds1003
 PIN vss.gds1004
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 15.318 31.922 15.518 ;
 END
 END vss.gds1004
 PIN vss.gds1005
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 15.278 30.95 15.478 ;
 END
 END vss.gds1005
 PIN vss.gds1006
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.314 13.152 30.37 13.352 ;
 END
 END vss.gds1006
 PIN vss.gds1007
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 13.14 32.214 13.34 ;
 END
 END vss.gds1007
 PIN vss.gds1008
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 13.0585 34.046 13.2585 ;
 END
 END vss.gds1008
 PIN vss.gds1009
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 13.0995 30.71 13.2995 ;
 END
 END vss.gds1009
 PIN vss.gds1010
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 14.773 33.198 14.973 ;
 END
 END vss.gds1010
 PIN vss.gds1011
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 13.513 33.198 13.713 ;
 END
 END vss.gds1011
 PIN vss.gds1012
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 14.018 30.95 14.218 ;
 END
 END vss.gds1012
 PIN vss.gds1013
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 10.993 33.198 11.193 ;
 END
 END vss.gds1013
 PIN vss.gds1014
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 12.253 33.198 12.453 ;
 END
 END vss.gds1014
 PIN vss.gds1015
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 13.14 32.894 13.34 ;
 END
 END vss.gds1015
 PIN vss.gds1016
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 12.758 30.95 12.958 ;
 END
 END vss.gds1016
 PIN vss.gds1017
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 12.9065 33.542 13.1065 ;
 END
 END vss.gds1017
 PIN vss.gds1018
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 13.14 31.55 13.34 ;
 END
 END vss.gds1018
 PIN vss.gds1019
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 13.152 33.866 13.352 ;
 END
 END vss.gds1019
 PIN vss.gds1020
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 13.0035 34.886 13.2035 ;
 END
 END vss.gds1020
 PIN vss.gds1021
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.49 13.1555 34.546 13.3555 ;
 END
 END vss.gds1021
 PIN vss.gds1022
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 12.996 32.47 13.196 ;
 END
 END vss.gds1022
 PIN vss.gds1023
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 13.0035 34.366 13.2035 ;
 END
 END vss.gds1023
 PIN vss.gds1024
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.038 12.883 35.078 13.083 ;
 END
 END vss.gds1024
 PIN vss.gds1025
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 32.648 13.18 32.704 13.38 ;
 RECT 32.9 13.183 32.956 13.383 ;
 RECT 33.572 14.216 33.628 14.369 ;
 RECT 31.052 14.196 31.108 14.369 ;
 RECT 31.22 14.169 31.276 14.369 ;
 RECT 32.816 14.213 32.872 14.378 ;
 RECT 32.648 14.213 32.704 14.378 ;
 RECT 31.892 14.213 31.948 14.378 ;
 RECT 31.724 14.213 31.78 14.378 ;
 RECT 33.572 11.696 33.628 11.849 ;
 RECT 31.052 11.676 31.108 11.849 ;
 RECT 31.22 11.649 31.276 11.849 ;
 RECT 32.816 11.693 32.872 11.858 ;
 RECT 32.648 11.693 32.704 11.858 ;
 RECT 31.892 11.693 31.948 11.858 ;
 RECT 31.724 11.693 31.78 11.858 ;
 RECT 33.572 12.956 33.628 13.109 ;
 RECT 31.052 12.936 31.108 13.109 ;
 RECT 31.22 12.909 31.276 13.109 ;
 RECT 32.816 12.953 32.872 13.118 ;
 RECT 32.648 12.953 32.704 13.118 ;
 RECT 31.892 12.953 31.948 13.118 ;
 RECT 31.724 12.953 31.78 13.118 ;
 RECT 33.572 15.476 33.628 15.629 ;
 RECT 31.052 15.456 31.108 15.629 ;
 RECT 31.22 15.429 31.276 15.629 ;
 RECT 32.816 15.473 32.872 15.638 ;
 RECT 32.648 15.473 32.704 15.638 ;
 RECT 31.892 15.473 31.948 15.638 ;
 RECT 31.724 15.473 31.78 15.638 ;
 RECT 32.648 10.66 32.704 10.86 ;
 RECT 32.9 10.663 32.956 10.863 ;
 RECT 32.648 11.92 32.704 12.12 ;
 RECT 32.9 11.923 32.956 12.123 ;
 RECT 32.648 14.44 32.704 14.64 ;
 RECT 32.9 14.443 32.956 14.643 ;
 RECT 31.388 13.529 31.444 13.729 ;
 RECT 31.22 13.529 31.276 13.729 ;
 RECT 32.06 13.739 32.116 13.939 ;
 RECT 32.48 13.739 32.536 13.939 ;
 RECT 33.908 14.8475 33.964 15.0475 ;
 RECT 33.404 15.0995 33.46 15.2995 ;
 RECT 32.06 14.999 32.116 15.199 ;
 RECT 32.48 14.999 32.536 15.199 ;
 RECT 31.388 14.789 31.444 14.989 ;
 RECT 31.22 14.789 31.276 14.989 ;
 RECT 30.716 14.923 30.772 15.123 ;
 RECT 31.388 12.269 31.444 12.469 ;
 RECT 31.22 12.269 31.276 12.469 ;
 RECT 32.06 12.479 32.116 12.679 ;
 RECT 32.48 12.479 32.536 12.679 ;
 RECT 30.716 12.403 30.772 12.603 ;
 RECT 33.404 12.5795 33.46 12.7795 ;
 RECT 33.908 12.3275 33.964 12.5275 ;
 RECT 33.404 11.3195 33.46 11.5195 ;
 RECT 33.908 11.0675 33.964 11.2675 ;
 RECT 31.388 11.009 31.444 11.209 ;
 RECT 31.22 11.009 31.276 11.209 ;
 RECT 30.716 11.143 30.772 11.343 ;
 RECT 32.06 11.219 32.116 11.419 ;
 RECT 32.48 11.219 32.536 11.419 ;
 RECT 30.716 13.663 30.772 13.863 ;
 RECT 33.404 13.8395 33.46 14.0395 ;
 RECT 33.908 13.5875 33.964 13.7875 ;
 RECT 30.548 12.975 30.604 13.175 ;
 RECT 30.38 12.913 30.436 13.113 ;
 RECT 32.228 13.1795 32.284 13.3795 ;
 RECT 34.916 12.994 34.972 13.194 ;
 RECT 34.748 13.0015 34.804 13.2015 ;
 RECT 34.58 12.994 34.636 13.194 ;
 RECT 34.412 12.994 34.468 13.194 ;
 RECT 34.244 12.994 34.3 13.194 ;
 RECT 35.084 12.994 35.14 13.194 ;
 RECT 34.076 13.109 34.132 13.309 ;
 END
 END vss.gds1025
 PIN vss.gds1026
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.122 13.0995 40.182 13.2995 ;
 END
 END vss.gds1026
 PIN vss.gds1027
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.754 13.0995 35.814 13.2995 ;
 END
 END vss.gds1027
 PIN vss.gds1028
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.09 13.0995 36.15 13.2995 ;
 END
 END vss.gds1028
 PIN vss.gds1029
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.258 13.0995 36.318 13.2995 ;
 END
 END vss.gds1029
 PIN vss.gds1030
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.426 13.0995 36.486 13.2995 ;
 END
 END vss.gds1030
 PIN vss.gds1031
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.762 13.0995 36.822 13.2995 ;
 END
 END vss.gds1031
 PIN vss.gds1032
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.93 13.0995 36.99 13.2995 ;
 END
 END vss.gds1032
 PIN vss.gds1033
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.098 13.0995 37.158 13.2995 ;
 END
 END vss.gds1033
 PIN vss.gds1034
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.434 13.0995 37.494 13.2995 ;
 END
 END vss.gds1034
 PIN vss.gds1035
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.602 13.0995 37.662 13.2995 ;
 END
 END vss.gds1035
 PIN vss.gds1036
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.77 13.0995 37.83 13.2995 ;
 END
 END vss.gds1036
 PIN vss.gds1037
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.106 13.0995 38.166 13.2995 ;
 END
 END vss.gds1037
 PIN vss.gds1038
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.274 13.0995 38.334 13.2995 ;
 END
 END vss.gds1038
 PIN vss.gds1039
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 13.0995 36.654 13.2995 ;
 END
 END vss.gds1039
 PIN vss.gds1040
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 13.0995 37.326 13.2995 ;
 END
 END vss.gds1040
 PIN vss.gds1041
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 13.0995 37.998 13.2995 ;
 END
 END vss.gds1041
 PIN vss.gds1042
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.442 13.0995 38.502 13.2995 ;
 END
 END vss.gds1042
 PIN vss.gds1043
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 13.0995 38.67 13.2995 ;
 END
 END vss.gds1043
 PIN vss.gds1044
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.778 13.0995 38.838 13.2995 ;
 END
 END vss.gds1044
 PIN vss.gds1045
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 13.0995 35.982 13.2995 ;
 END
 END vss.gds1045
 PIN vss.gds1046
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.946 13.0995 39.006 13.2995 ;
 END
 END vss.gds1046
 PIN vss.gds1047
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.586 13.0995 35.646 13.2995 ;
 END
 END vss.gds1047
 PIN vss.gds1048
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.45 13.0995 39.51 13.2995 ;
 END
 END vss.gds1048
 PIN vss.gds1049
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.618 13.0995 39.678 13.2995 ;
 END
 END vss.gds1049
 PIN vss.gds1050
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.114 13.0995 39.174 13.2995 ;
 END
 END vss.gds1050
 PIN vss.gds1051
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.786 13.0995 39.846 13.2995 ;
 END
 END vss.gds1051
 PIN vss.gds1052
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 13.0995 40.014 13.2995 ;
 END
 END vss.gds1052
 PIN vss.gds1053
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.418 13.0995 35.478 13.2995 ;
 END
 END vss.gds1053
 PIN vss.gds1054
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 13.021 35.31 13.221 ;
 END
 END vss.gds1054
 PIN vss.gds1055
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 13.0995 39.342 13.2995 ;
 END
 END vss.gds1055
 PIN vss.gds1056
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.91 13.0995 44.97 13.2995 ;
 END
 END vss.gds1056
 PIN vss.gds1057
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.742 13.0995 44.802 13.2995 ;
 END
 END vss.gds1057
 PIN vss.gds1058
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.574 13.0995 44.634 13.2995 ;
 END
 END vss.gds1058
 PIN vss.gds1059
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.238 13.0995 44.298 13.2995 ;
 END
 END vss.gds1059
 PIN vss.gds1060
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.07 13.0995 44.13 13.2995 ;
 END
 END vss.gds1060
 PIN vss.gds1061
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.902 13.0995 43.962 13.2995 ;
 END
 END vss.gds1061
 PIN vss.gds1062
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.566 13.0995 43.626 13.2995 ;
 END
 END vss.gds1062
 PIN vss.gds1063
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.398 13.0995 43.458 13.2995 ;
 END
 END vss.gds1063
 PIN vss.gds1064
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.23 13.0995 43.29 13.2995 ;
 END
 END vss.gds1064
 PIN vss.gds1065
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.894 13.0995 42.954 13.2995 ;
 END
 END vss.gds1065
 PIN vss.gds1066
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.726 13.0995 42.786 13.2995 ;
 END
 END vss.gds1066
 PIN vss.gds1067
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.558 13.0995 42.618 13.2995 ;
 END
 END vss.gds1067
 PIN vss.gds1068
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.222 13.0995 42.282 13.2995 ;
 END
 END vss.gds1068
 PIN vss.gds1069
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.054 13.0995 42.114 13.2995 ;
 END
 END vss.gds1069
 PIN vss.gds1070
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.886 13.0995 41.946 13.2995 ;
 END
 END vss.gds1070
 PIN vss.gds1071
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.55 13.0995 41.61 13.2995 ;
 END
 END vss.gds1071
 PIN vss.gds1072
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.382 13.0995 41.442 13.2995 ;
 END
 END vss.gds1072
 PIN vss.gds1073
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.214 13.0995 41.274 13.2995 ;
 END
 END vss.gds1073
 PIN vss.gds1074
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.29 13.0995 40.35 13.2995 ;
 END
 END vss.gds1074
 PIN vss.gds1075
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.458 13.0995 40.518 13.2995 ;
 END
 END vss.gds1075
 PIN vss.gds1076
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 13.0995 45.138 13.2995 ;
 END
 END vss.gds1076
 PIN vss.gds1077
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 13.0995 44.466 13.2995 ;
 END
 END vss.gds1077
 PIN vss.gds1078
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 13.0995 43.794 13.2995 ;
 END
 END vss.gds1078
 PIN vss.gds1079
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 13.0995 43.122 13.2995 ;
 END
 END vss.gds1079
 PIN vss.gds1080
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 13.0995 42.45 13.2995 ;
 END
 END vss.gds1080
 PIN vss.gds1081
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 13.0995 41.778 13.2995 ;
 END
 END vss.gds1081
 PIN vss.gds1082
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 13.0995 40.686 13.2995 ;
 END
 END vss.gds1082
 PIN vss.gds1083
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 40.964 13.676 41.02 13.876 ;
 RECT 40.964 14.936 41.02 15.136 ;
 RECT 40.964 12.416 41.02 12.616 ;
 RECT 40.964 11.156 41.02 11.356 ;
 RECT 40.796 13.046 40.852 13.246 ;
 END
 END vss.gds1083
 PIN vss.gds1084
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 12.798 48.974 12.998 ;
 END
 END vss.gds1084
 PIN vss.gds1085
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 11.498 48.002 11.698 ;
 END
 END vss.gds1085
 PIN vss.gds1086
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 11.538 48.974 11.738 ;
 END
 END vss.gds1086
 PIN vss.gds1087
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 14.058 48.974 14.258 ;
 END
 END vss.gds1087
 PIN vss.gds1088
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 15.318 48.974 15.518 ;
 END
 END vss.gds1088
 PIN vss.gds1089
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 15.278 48.002 15.478 ;
 END
 END vss.gds1089
 PIN vss.gds1090
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.366 13.152 47.422 13.352 ;
 END
 END vss.gds1090
 PIN vss.gds1091
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.254 13.0995 46.314 13.2995 ;
 END
 END vss.gds1091
 PIN vss.gds1092
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.086 13.0995 46.146 13.2995 ;
 END
 END vss.gds1092
 PIN vss.gds1093
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.918 13.0995 45.978 13.2995 ;
 END
 END vss.gds1093
 PIN vss.gds1094
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.582 13.0995 45.642 13.2995 ;
 END
 END vss.gds1094
 PIN vss.gds1095
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.414 13.0995 45.474 13.2995 ;
 END
 END vss.gds1095
 PIN vss.gds1096
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.246 13.0995 45.306 13.2995 ;
 END
 END vss.gds1096
 PIN vss.gds1097
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 13.1555 47.162 13.3555 ;
 END
 END vss.gds1097
 PIN vss.gds1098
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 13.021 46.482 13.221 ;
 END
 END vss.gds1098
 PIN vss.gds1099
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 13.0995 45.81 13.2995 ;
 END
 END vss.gds1099
 PIN vss.gds1100
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 13.0035 46.922 13.2035 ;
 END
 END vss.gds1100
 PIN vss.gds1101
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 12.883 46.694 13.083 ;
 END
 END vss.gds1101
 PIN vss.gds1102
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 13.0995 47.762 13.2995 ;
 END
 END vss.gds1102
 PIN vss.gds1103
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 13.14 49.266 13.34 ;
 END
 END vss.gds1103
 PIN vss.gds1104
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 13.14 48.602 13.34 ;
 END
 END vss.gds1104
 PIN vss.gds1105
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 14.773 50.25 14.973 ;
 END
 END vss.gds1105
 PIN vss.gds1106
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 13.513 50.25 13.713 ;
 END
 END vss.gds1106
 PIN vss.gds1107
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 12.253 50.25 12.453 ;
 END
 END vss.gds1107
 PIN vss.gds1108
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 14.018 48.002 14.218 ;
 END
 END vss.gds1108
 PIN vss.gds1109
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 13.14 49.946 13.34 ;
 END
 END vss.gds1109
 PIN vss.gds1110
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 12.758 48.002 12.958 ;
 END
 END vss.gds1110
 PIN vss.gds1111
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 10.993 50.25 11.193 ;
 END
 END vss.gds1111
 PIN vss.gds1112
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 12.996 49.522 13.196 ;
 END
 END vss.gds1112
 PIN vss.gds1113
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 49.7 13.18 49.756 13.38 ;
 RECT 49.952 13.183 50.008 13.383 ;
 RECT 48.104 14.196 48.16 14.369 ;
 RECT 48.272 14.169 48.328 14.369 ;
 RECT 49.868 14.213 49.924 14.378 ;
 RECT 49.7 14.213 49.756 14.378 ;
 RECT 48.944 14.213 49 14.378 ;
 RECT 48.776 14.213 48.832 14.378 ;
 RECT 48.104 11.676 48.16 11.849 ;
 RECT 48.272 11.649 48.328 11.849 ;
 RECT 49.868 11.693 49.924 11.858 ;
 RECT 49.7 11.693 49.756 11.858 ;
 RECT 48.944 11.693 49 11.858 ;
 RECT 48.776 11.693 48.832 11.858 ;
 RECT 48.104 12.936 48.16 13.109 ;
 RECT 48.272 12.909 48.328 13.109 ;
 RECT 49.868 12.953 49.924 13.118 ;
 RECT 49.7 12.953 49.756 13.118 ;
 RECT 48.944 12.953 49 13.118 ;
 RECT 48.776 12.953 48.832 13.118 ;
 RECT 48.104 15.456 48.16 15.629 ;
 RECT 48.272 15.429 48.328 15.629 ;
 RECT 49.868 15.473 49.924 15.638 ;
 RECT 49.7 15.473 49.756 15.638 ;
 RECT 48.944 15.473 49 15.638 ;
 RECT 48.776 15.473 48.832 15.638 ;
 RECT 49.7 10.66 49.756 10.86 ;
 RECT 49.952 10.663 50.008 10.863 ;
 RECT 48.44 11.009 48.496 11.209 ;
 RECT 48.272 11.009 48.328 11.209 ;
 RECT 49.7 11.92 49.756 12.12 ;
 RECT 49.952 11.923 50.008 12.123 ;
 RECT 49.7 14.44 49.756 14.64 ;
 RECT 49.952 14.443 50.008 14.643 ;
 RECT 48.44 13.529 48.496 13.729 ;
 RECT 48.272 13.529 48.328 13.729 ;
 RECT 49.112 13.739 49.168 13.939 ;
 RECT 49.532 13.739 49.588 13.939 ;
 RECT 48.44 12.269 48.496 12.469 ;
 RECT 48.272 12.269 48.328 12.469 ;
 RECT 49.112 12.479 49.168 12.679 ;
 RECT 49.532 12.479 49.588 12.679 ;
 RECT 49.112 14.999 49.168 15.199 ;
 RECT 49.532 14.999 49.588 15.199 ;
 RECT 48.44 14.789 48.496 14.989 ;
 RECT 48.272 14.789 48.328 14.989 ;
 RECT 47.768 14.923 47.824 15.123 ;
 RECT 47.768 12.403 47.824 12.603 ;
 RECT 47.768 11.143 47.824 11.343 ;
 RECT 49.112 11.219 49.168 11.419 ;
 RECT 49.532 11.219 49.588 11.419 ;
 RECT 47.768 13.663 47.824 13.863 ;
 RECT 47.6 12.975 47.656 13.175 ;
 RECT 47.432 12.913 47.488 13.113 ;
 RECT 47.264 12.964 47.32 13.164 ;
 RECT 46.928 12.964 46.984 13.164 ;
 RECT 47.096 12.964 47.152 13.164 ;
 RECT 49.28 13.1795 49.336 13.3795 ;
 RECT 46.592 12.994 46.648 13.194 ;
 RECT 46.76 12.994 46.816 13.194 ;
 END
 END vss.gds1113
 PIN vss.gds1114
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.638 13.0995 52.698 13.2995 ;
 END
 END vss.gds1114
 PIN vss.gds1115
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.806 13.0995 52.866 13.2995 ;
 END
 END vss.gds1115
 PIN vss.gds1116
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.142 13.0995 53.202 13.2995 ;
 END
 END vss.gds1116
 PIN vss.gds1117
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.31 13.0995 53.37 13.2995 ;
 END
 END vss.gds1117
 PIN vss.gds1118
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.478 13.0995 53.538 13.2995 ;
 END
 END vss.gds1118
 PIN vss.gds1119
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.814 13.0995 53.874 13.2995 ;
 END
 END vss.gds1119
 PIN vss.gds1120
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.982 13.0995 54.042 13.2995 ;
 END
 END vss.gds1120
 PIN vss.gds1121
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.15 13.0995 54.21 13.2995 ;
 END
 END vss.gds1121
 PIN vss.gds1122
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.486 13.0995 54.546 13.2995 ;
 END
 END vss.gds1122
 PIN vss.gds1123
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.654 13.0995 54.714 13.2995 ;
 END
 END vss.gds1123
 PIN vss.gds1124
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.822 13.0995 54.882 13.2995 ;
 END
 END vss.gds1124
 PIN vss.gds1125
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.158 13.0995 55.218 13.2995 ;
 END
 END vss.gds1125
 PIN vss.gds1126
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 13.0995 55.05 13.2995 ;
 END
 END vss.gds1126
 PIN vss.gds1127
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 13.0995 54.378 13.2995 ;
 END
 END vss.gds1127
 PIN vss.gds1128
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 13.152 50.918 13.352 ;
 END
 END vss.gds1128
 PIN vss.gds1129
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 13.0995 53.706 13.2995 ;
 END
 END vss.gds1129
 PIN vss.gds1130
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 13.0585 51.098 13.2585 ;
 END
 END vss.gds1130
 PIN vss.gds1131
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 13.0995 53.034 13.2995 ;
 END
 END vss.gds1131
 PIN vss.gds1132
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 13.0035 51.938 13.2035 ;
 END
 END vss.gds1132
 PIN vss.gds1133
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.542 13.1555 51.598 13.3555 ;
 END
 END vss.gds1133
 PIN vss.gds1134
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 13.0035 51.418 13.2035 ;
 END
 END vss.gds1134
 PIN vss.gds1135
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 12.9065 50.594 13.1065 ;
 END
 END vss.gds1135
 PIN vss.gds1136
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.09 12.883 52.13 13.083 ;
 END
 END vss.gds1136
 PIN vss.gds1137
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.47 13.0995 52.53 13.2995 ;
 END
 END vss.gds1137
 PIN vss.gds1138
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 13.021 52.362 13.221 ;
 END
 END vss.gds1138
 PIN vss.gds1139
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 50.624 14.216 50.68 14.369 ;
 RECT 50.624 11.696 50.68 11.849 ;
 RECT 50.624 12.956 50.68 13.109 ;
 RECT 50.624 15.476 50.68 15.629 ;
 RECT 50.96 14.8475 51.016 15.0475 ;
 RECT 50.456 15.0995 50.512 15.2995 ;
 RECT 50.456 12.5795 50.512 12.7795 ;
 RECT 50.96 12.3275 51.016 12.5275 ;
 RECT 50.456 13.8395 50.512 14.0395 ;
 RECT 50.96 13.5875 51.016 13.7875 ;
 RECT 50.456 11.3195 50.512 11.5195 ;
 RECT 50.96 11.0675 51.016 11.2675 ;
 RECT 51.968 12.994 52.024 13.194 ;
 RECT 51.8 13.0015 51.856 13.2015 ;
 RECT 51.632 12.994 51.688 13.194 ;
 RECT 51.464 12.994 51.52 13.194 ;
 RECT 51.296 12.994 51.352 13.194 ;
 RECT 52.136 12.994 52.192 13.194 ;
 RECT 51.128 13.109 51.184 13.309 ;
 END
 END vss.gds1139
 PIN vss.gds1140
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.946 13.0995 60.006 13.2995 ;
 END
 END vss.gds1140
 PIN vss.gds1141
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.778 13.0995 59.838 13.2995 ;
 END
 END vss.gds1141
 PIN vss.gds1142
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.61 13.0995 59.67 13.2995 ;
 END
 END vss.gds1142
 PIN vss.gds1143
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.274 13.0995 59.334 13.2995 ;
 END
 END vss.gds1143
 PIN vss.gds1144
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.106 13.0995 59.166 13.2995 ;
 END
 END vss.gds1144
 PIN vss.gds1145
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.938 13.0995 58.998 13.2995 ;
 END
 END vss.gds1145
 PIN vss.gds1146
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.602 13.0995 58.662 13.2995 ;
 END
 END vss.gds1146
 PIN vss.gds1147
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.434 13.0995 58.494 13.2995 ;
 END
 END vss.gds1147
 PIN vss.gds1148
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.266 13.0995 58.326 13.2995 ;
 END
 END vss.gds1148
 PIN vss.gds1149
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.326 13.0995 55.386 13.2995 ;
 END
 END vss.gds1149
 PIN vss.gds1150
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.494 13.0995 55.554 13.2995 ;
 END
 END vss.gds1150
 PIN vss.gds1151
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 13.0995 60.174 13.2995 ;
 END
 END vss.gds1151
 PIN vss.gds1152
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 13.0995 59.502 13.2995 ;
 END
 END vss.gds1152
 PIN vss.gds1153
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 13.0995 58.83 13.2995 ;
 END
 END vss.gds1153
 PIN vss.gds1154
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 13.0995 55.722 13.2995 ;
 END
 END vss.gds1154
 PIN vss.gds1155
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.83 13.0995 55.89 13.2995 ;
 END
 END vss.gds1155
 PIN vss.gds1156
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.998 13.0995 56.058 13.2995 ;
 END
 END vss.gds1156
 PIN vss.gds1157
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.166 13.0995 56.226 13.2995 ;
 END
 END vss.gds1157
 PIN vss.gds1158
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 13.0995 56.394 13.2995 ;
 END
 END vss.gds1158
 PIN vss.gds1159
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.502 13.0995 56.562 13.2995 ;
 END
 END vss.gds1159
 PIN vss.gds1160
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.67 13.0995 56.73 13.2995 ;
 END
 END vss.gds1160
 PIN vss.gds1161
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.838 13.0995 56.898 13.2995 ;
 END
 END vss.gds1161
 PIN vss.gds1162
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.342 13.0995 57.402 13.2995 ;
 END
 END vss.gds1162
 PIN vss.gds1163
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.51 13.0995 57.57 13.2995 ;
 END
 END vss.gds1163
 PIN vss.gds1164
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 13.0995 57.738 13.2995 ;
 END
 END vss.gds1164
 PIN vss.gds1165
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.174 13.0995 57.234 13.2995 ;
 END
 END vss.gds1165
 PIN vss.gds1166
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 13.0995 57.066 13.2995 ;
 END
 END vss.gds1166
 PIN vss.gds1167
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 58.016 13.676 58.072 13.876 ;
 RECT 58.016 12.416 58.072 12.616 ;
 RECT 58.016 14.936 58.072 15.136 ;
 RECT 58.016 11.156 58.072 11.356 ;
 RECT 57.848 13.046 57.904 13.246 ;
 END
 END vss.gds1167
 PIN vss.gds1168
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 11.498 65.054 11.698 ;
 END
 END vss.gds1168
 PIN vss.gds1169
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 14.018 65.054 14.218 ;
 END
 END vss.gds1169
 PIN vss.gds1170
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 15.278 65.054 15.478 ;
 END
 END vss.gds1170
 PIN vss.gds1171
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 13.1555 64.214 13.3555 ;
 END
 END vss.gds1171
 PIN vss.gds1172
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.418 13.152 64.474 13.352 ;
 END
 END vss.gds1172
 PIN vss.gds1173
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.306 13.0995 63.366 13.2995 ;
 END
 END vss.gds1173
 PIN vss.gds1174
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.138 13.0995 63.198 13.2995 ;
 END
 END vss.gds1174
 PIN vss.gds1175
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.97 13.0995 63.03 13.2995 ;
 END
 END vss.gds1175
 PIN vss.gds1176
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.634 13.0995 62.694 13.2995 ;
 END
 END vss.gds1176
 PIN vss.gds1177
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.466 13.0995 62.526 13.2995 ;
 END
 END vss.gds1177
 PIN vss.gds1178
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.298 13.0995 62.358 13.2995 ;
 END
 END vss.gds1178
 PIN vss.gds1179
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.962 13.0995 62.022 13.2995 ;
 END
 END vss.gds1179
 PIN vss.gds1180
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.794 13.0995 61.854 13.2995 ;
 END
 END vss.gds1180
 PIN vss.gds1181
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.626 13.0995 61.686 13.2995 ;
 END
 END vss.gds1181
 PIN vss.gds1182
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.29 13.0995 61.35 13.2995 ;
 END
 END vss.gds1182
 PIN vss.gds1183
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.122 13.0995 61.182 13.2995 ;
 END
 END vss.gds1183
 PIN vss.gds1184
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.954 13.0995 61.014 13.2995 ;
 END
 END vss.gds1184
 PIN vss.gds1185
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.618 13.0995 60.678 13.2995 ;
 END
 END vss.gds1185
 PIN vss.gds1186
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.45 13.0995 60.51 13.2995 ;
 END
 END vss.gds1186
 PIN vss.gds1187
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.282 13.0995 60.342 13.2995 ;
 END
 END vss.gds1187
 PIN vss.gds1188
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 13.021 63.534 13.221 ;
 END
 END vss.gds1188
 PIN vss.gds1189
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 13.0995 62.862 13.2995 ;
 END
 END vss.gds1189
 PIN vss.gds1190
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 13.0995 62.19 13.2995 ;
 END
 END vss.gds1190
 PIN vss.gds1191
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 13.0995 61.518 13.2995 ;
 END
 END vss.gds1191
 PIN vss.gds1192
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 13.0995 60.846 13.2995 ;
 END
 END vss.gds1192
 PIN vss.gds1193
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 13.0035 63.974 13.2035 ;
 END
 END vss.gds1193
 PIN vss.gds1194
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 12.883 63.746 13.083 ;
 END
 END vss.gds1194
 PIN vss.gds1195
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 13.0995 64.814 13.2995 ;
 END
 END vss.gds1195
 PIN vss.gds1196
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 12.758 65.054 12.958 ;
 END
 END vss.gds1196
 PIN vss.gds1197
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 65.156 14.196 65.212 14.369 ;
 RECT 65.156 11.676 65.212 11.849 ;
 RECT 65.156 12.936 65.212 13.109 ;
 RECT 65.156 15.456 65.212 15.629 ;
 RECT 64.82 14.923 64.876 15.123 ;
 RECT 64.82 13.663 64.876 13.863 ;
 RECT 64.82 12.403 64.876 12.603 ;
 RECT 64.82 11.143 64.876 11.343 ;
 RECT 64.652 12.975 64.708 13.175 ;
 RECT 64.484 12.913 64.54 13.113 ;
 RECT 64.316 12.964 64.372 13.164 ;
 RECT 64.148 12.964 64.204 13.164 ;
 RECT 63.98 12.964 64.036 13.164 ;
 RECT 63.644 12.994 63.7 13.194 ;
 RECT 63.812 12.994 63.868 13.194 ;
 END
 END vss.gds1197
 PIN vss.gds1198
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 12.798 66.026 12.998 ;
 END
 END vss.gds1198
 PIN vss.gds1199
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 11.538 66.026 11.738 ;
 END
 END vss.gds1199
 PIN vss.gds1200
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 14.058 66.026 14.258 ;
 END
 END vss.gds1200
 PIN vss.gds1201
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 15.318 66.026 15.518 ;
 END
 END vss.gds1201
 PIN vss.gds1202
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.69 13.0995 69.75 13.2995 ;
 END
 END vss.gds1202
 PIN vss.gds1203
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.858 13.0995 69.918 13.2995 ;
 END
 END vss.gds1203
 PIN vss.gds1204
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.194 13.0995 70.254 13.2995 ;
 END
 END vss.gds1204
 PIN vss.gds1205
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 13.0585 68.15 13.2585 ;
 END
 END vss.gds1205
 PIN vss.gds1206
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 13.14 66.318 13.34 ;
 END
 END vss.gds1206
 PIN vss.gds1207
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 13.0995 70.086 13.2995 ;
 END
 END vss.gds1207
 PIN vss.gds1208
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 13.14 66.998 13.34 ;
 END
 END vss.gds1208
 PIN vss.gds1209
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 14.773 67.302 14.973 ;
 END
 END vss.gds1209
 PIN vss.gds1210
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 13.513 67.302 13.713 ;
 END
 END vss.gds1210
 PIN vss.gds1211
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 12.253 67.302 12.453 ;
 END
 END vss.gds1211
 PIN vss.gds1212
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 10.993 67.302 11.193 ;
 END
 END vss.gds1212
 PIN vss.gds1213
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 13.14 65.654 13.34 ;
 END
 END vss.gds1213
 PIN vss.gds1214
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 12.9065 67.646 13.1065 ;
 END
 END vss.gds1214
 PIN vss.gds1215
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 12.996 66.574 13.196 ;
 END
 END vss.gds1215
 PIN vss.gds1216
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 13.152 67.97 13.352 ;
 END
 END vss.gds1216
 PIN vss.gds1217
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 13.0035 68.99 13.2035 ;
 END
 END vss.gds1217
 PIN vss.gds1218
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.594 13.1555 68.65 13.3555 ;
 END
 END vss.gds1218
 PIN vss.gds1219
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 13.0035 68.47 13.2035 ;
 END
 END vss.gds1219
 PIN vss.gds1220
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.142 12.883 69.182 13.083 ;
 END
 END vss.gds1220
 PIN vss.gds1221
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.522 13.0995 69.582 13.2995 ;
 END
 END vss.gds1221
 PIN vss.gds1222
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 13.021 69.414 13.221 ;
 END
 END vss.gds1222
 PIN vss.gds1223
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 66.752 10.66 66.808 10.86 ;
 RECT 67.004 10.663 67.06 10.863 ;
 RECT 66.752 13.18 66.808 13.38 ;
 RECT 67.004 13.183 67.06 13.383 ;
 RECT 67.676 14.216 67.732 14.369 ;
 RECT 65.324 14.169 65.38 14.369 ;
 RECT 66.92 14.213 66.976 14.378 ;
 RECT 66.752 14.213 66.808 14.378 ;
 RECT 65.996 14.213 66.052 14.378 ;
 RECT 65.828 14.213 65.884 14.378 ;
 RECT 67.676 11.696 67.732 11.849 ;
 RECT 65.324 11.649 65.38 11.849 ;
 RECT 66.92 11.693 66.976 11.858 ;
 RECT 66.752 11.693 66.808 11.858 ;
 RECT 65.996 11.693 66.052 11.858 ;
 RECT 65.828 11.693 65.884 11.858 ;
 RECT 67.676 12.956 67.732 13.109 ;
 RECT 65.324 12.909 65.38 13.109 ;
 RECT 66.92 12.953 66.976 13.118 ;
 RECT 66.752 12.953 66.808 13.118 ;
 RECT 65.996 12.953 66.052 13.118 ;
 RECT 65.828 12.953 65.884 13.118 ;
 RECT 67.676 15.476 67.732 15.629 ;
 RECT 65.324 15.429 65.38 15.629 ;
 RECT 66.92 15.473 66.976 15.638 ;
 RECT 66.752 15.473 66.808 15.638 ;
 RECT 65.996 15.473 66.052 15.638 ;
 RECT 65.828 15.473 65.884 15.638 ;
 RECT 66.752 11.92 66.808 12.12 ;
 RECT 67.004 11.923 67.06 12.123 ;
 RECT 66.752 14.44 66.808 14.64 ;
 RECT 67.004 14.443 67.06 14.643 ;
 RECT 65.492 13.529 65.548 13.729 ;
 RECT 65.324 13.529 65.38 13.729 ;
 RECT 67.508 13.8395 67.564 14.0395 ;
 RECT 68.012 13.5875 68.068 13.7875 ;
 RECT 68.012 14.8475 68.068 15.0475 ;
 RECT 67.508 15.0995 67.564 15.2995 ;
 RECT 66.164 14.999 66.22 15.199 ;
 RECT 66.584 14.999 66.64 15.199 ;
 RECT 65.492 14.789 65.548 14.989 ;
 RECT 65.324 14.789 65.38 14.989 ;
 RECT 66.164 13.739 66.22 13.939 ;
 RECT 66.584 13.739 66.64 13.939 ;
 RECT 65.492 12.269 65.548 12.469 ;
 RECT 65.324 12.269 65.38 12.469 ;
 RECT 66.164 12.479 66.22 12.679 ;
 RECT 66.584 12.479 66.64 12.679 ;
 RECT 67.508 12.5795 67.564 12.7795 ;
 RECT 68.012 12.3275 68.068 12.5275 ;
 RECT 68.012 11.0675 68.068 11.2675 ;
 RECT 67.508 11.3195 67.564 11.5195 ;
 RECT 66.164 11.219 66.22 11.419 ;
 RECT 66.584 11.219 66.64 11.419 ;
 RECT 65.492 11.009 65.548 11.209 ;
 RECT 65.324 11.009 65.38 11.209 ;
 RECT 66.332 13.1795 66.388 13.3795 ;
 RECT 69.02 12.994 69.076 13.194 ;
 RECT 68.852 13.0015 68.908 13.2015 ;
 RECT 68.684 12.994 68.74 13.194 ;
 RECT 68.516 12.994 68.572 13.194 ;
 RECT 68.348 12.994 68.404 13.194 ;
 RECT 69.188 12.994 69.244 13.194 ;
 RECT 68.18 13.109 68.236 13.309 ;
 END
 END vss.gds1223
 PIN vss.gds1224
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.362 13.0995 70.422 13.2995 ;
 END
 END vss.gds1224
 PIN vss.gds1225
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.53 13.0995 70.59 13.2995 ;
 END
 END vss.gds1225
 PIN vss.gds1226
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.866 13.0995 70.926 13.2995 ;
 END
 END vss.gds1226
 PIN vss.gds1227
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.034 13.0995 71.094 13.2995 ;
 END
 END vss.gds1227
 PIN vss.gds1228
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.202 13.0995 71.262 13.2995 ;
 END
 END vss.gds1228
 PIN vss.gds1229
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.538 13.0995 71.598 13.2995 ;
 END
 END vss.gds1229
 PIN vss.gds1230
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.706 13.0995 71.766 13.2995 ;
 END
 END vss.gds1230
 PIN vss.gds1231
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.874 13.0995 71.934 13.2995 ;
 END
 END vss.gds1231
 PIN vss.gds1232
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.21 13.0995 72.27 13.2995 ;
 END
 END vss.gds1232
 PIN vss.gds1233
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.378 13.0995 72.438 13.2995 ;
 END
 END vss.gds1233
 PIN vss.gds1234
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.546 13.0995 72.606 13.2995 ;
 END
 END vss.gds1234
 PIN vss.gds1235
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.882 13.0995 72.942 13.2995 ;
 END
 END vss.gds1235
 PIN vss.gds1236
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.05 13.0995 73.11 13.2995 ;
 END
 END vss.gds1236
 PIN vss.gds1237
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 13.0995 71.43 13.2995 ;
 END
 END vss.gds1237
 PIN vss.gds1238
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 13.0995 72.102 13.2995 ;
 END
 END vss.gds1238
 PIN vss.gds1239
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 13.0995 72.774 13.2995 ;
 END
 END vss.gds1239
 PIN vss.gds1240
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 13.0995 70.758 13.2995 ;
 END
 END vss.gds1240
 PIN vss.gds1241
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.554 13.0995 73.614 13.2995 ;
 END
 END vss.gds1241
 PIN vss.gds1242
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.722 13.0995 73.782 13.2995 ;
 END
 END vss.gds1242
 PIN vss.gds1243
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 13.0995 73.446 13.2995 ;
 END
 END vss.gds1243
 PIN vss.gds1244
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.218 13.0995 73.278 13.2995 ;
 END
 END vss.gds1244
 PIN vss.gds1245
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.89 13.0995 73.95 13.2995 ;
 END
 END vss.gds1245
 PIN vss.gds1246
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.394 13.0995 74.454 13.2995 ;
 END
 END vss.gds1246
 PIN vss.gds1247
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 13.0995 74.118 13.2995 ;
 END
 END vss.gds1247
 PIN vss.gds1248
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.562 13.0995 74.622 13.2995 ;
 END
 END vss.gds1248
 PIN vss.gds1249
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 13.0995 74.79 13.2995 ;
 END
 END vss.gds1249
 PIN vss.gds1250
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.226 13.0995 74.286 13.2995 ;
 END
 END vss.gds1250
 PIN vss.gds1251
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 18.553 2.962 18.753 ;
 END
 END vss.gds1251
 PIN vss.gds1252
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 19.813 2.962 20.013 ;
 END
 END vss.gds1252
 PIN vss.gds1253
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 16.033 2.962 16.233 ;
 END
 END vss.gds1253
 PIN vss.gds1254
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 19.412 3.142 19.612 ;
 END
 END vss.gds1254
 PIN vss.gds1255
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 17.293 2.962 17.493 ;
 END
 END vss.gds1255
 PIN vss.gds1256
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 16.892 3.142 17.092 ;
 END
 END vss.gds1256
 PIN vss.gds1257
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 18.152 3.142 18.352 ;
 END
 END vss.gds1257
 PIN vss.gds1258
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 15.632 3.142 15.832 ;
 END
 END vss.gds1258
 PIN vss.gds1259
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 17.517 0.942 17.717 ;
 END
 END vss.gds1259
 PIN vss.gds1260
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.286 17.923 3.326 18.123 ;
 END
 END vss.gds1260
 PIN vss.gds1261
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 18.5015 4.194 18.7015 ;
 END
 END vss.gds1261
 PIN vss.gds1262
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 17.923 5.074 18.123 ;
 END
 END vss.gds1262
 PIN vss.gds1263
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 17.6175 0.718 17.8175 ;
 END
 END vss.gds1263
 PIN vss.gds1264
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.442 17.517 4.482 17.717 ;
 END
 END vss.gds1264
 PIN vss.gds1265
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.57 17.72 4.61 17.92 ;
 END
 END vss.gds1265
 PIN vss.gds1266
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 17.517 4.882 17.717 ;
 END
 END vss.gds1266
 PIN vss.gds1267
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 17.718 0.602 17.918 ;
 END
 END vss.gds1267
 PIN vss.gds1268
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 17.9465 2.122 18.1465 ;
 END
 END vss.gds1268
 PIN vss.gds1269
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 18.061 1.282 18.261 ;
 END
 END vss.gds1269
 PIN vss.gds1270
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 18.2955 1.462 18.4955 ;
 END
 END vss.gds1270
 PIN vss.gds1271
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.414 18.199 3.454 18.399 ;
 END
 END vss.gds1271
 PIN vss.gds1272
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.562 18.199 3.602 18.399 ;
 END
 END vss.gds1272
 PIN vss.gds1273
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 17.858 2.302 18.058 ;
 END
 END vss.gds1273
 PIN vss.gds1274
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 17.8195 4.002 18.0195 ;
 END
 END vss.gds1274
 PIN vss.gds1275
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 17.8195 5.282 18.0195 ;
 END
 END vss.gds1275
 PIN vss.gds1276
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 17.939 0.29 18.139 ;
 END
 END vss.gds1276
 PIN vss.gds1277
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.754 17.923 3.794 18.123 ;
 END
 END vss.gds1277
 PIN vss.gds1278
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 2.408 19.8135 2.464 20.0135 ;
 RECT 2.576 19.8135 2.632 20.0135 ;
 RECT 2.996 19.8135 3.052 20.0135 ;
 RECT 0.812 19.905 0.868 20.105 ;
 RECT 3.332 19.905 3.388 20.105 ;
 RECT 2.408 18.5535 2.464 18.7535 ;
 RECT 2.576 18.5535 2.632 18.7535 ;
 RECT 2.996 18.5535 3.052 18.7535 ;
 RECT 3.332 18.645 3.388 18.845 ;
 RECT 3.5 18.6015 3.556 18.8015 ;
 RECT 0.98 18.4685 1.036 18.6685 ;
 RECT 2.072 18.469 2.128 18.669 ;
 RECT 2.408 17.2935 2.464 17.4935 ;
 RECT 2.576 17.2935 2.632 17.4935 ;
 RECT 2.996 17.2935 3.052 17.4935 ;
 RECT 0.812 17.385 0.868 17.585 ;
 RECT 3.332 17.385 3.388 17.585 ;
 RECT 2.576 16.0335 2.632 16.2335 ;
 RECT 2.408 16.0335 2.464 16.2335 ;
 RECT 2.996 16.0335 3.052 16.2335 ;
 RECT 3.332 16.125 3.388 16.325 ;
 RECT 3.5 16.0815 3.556 16.2815 ;
 RECT 0.98 15.9485 1.036 16.1485 ;
 RECT 2.072 15.949 2.128 16.149 ;
 RECT 0.392 16.039 0.448 16.239 ;
 RECT 0.812 16.125 0.868 16.325 ;
 RECT 0.644 16.039 0.7 16.239 ;
 RECT 1.232 16.039 1.288 16.239 ;
 RECT 1.4 16.039 1.456 16.239 ;
 RECT 1.568 16.039 1.624 16.239 ;
 RECT 1.82 16.039 1.876 16.239 ;
 RECT 2.24 16.039 2.296 16.239 ;
 RECT 2.744 15.949 2.8 16.149 ;
 RECT 3.164 16.039 3.22 16.239 ;
 RECT 3.92 16.039 3.976 16.239 ;
 RECT 3.752 16.309 3.808 16.509 ;
 RECT 4.508 16.2385 4.564 16.4385 ;
 RECT 3.5 17.3415 3.556 17.5415 ;
 RECT 0.392 17.299 0.448 17.499 ;
 RECT 0.644 17.299 0.7 17.499 ;
 RECT 1.232 17.299 1.288 17.499 ;
 RECT 0.98 17.2085 1.036 17.4085 ;
 RECT 1.4 17.299 1.456 17.499 ;
 RECT 1.568 17.299 1.624 17.499 ;
 RECT 2.072 17.209 2.128 17.409 ;
 RECT 1.82 17.299 1.876 17.499 ;
 RECT 2.744 17.209 2.8 17.409 ;
 RECT 3.164 17.299 3.22 17.499 ;
 RECT 3.92 17.299 3.976 17.499 ;
 RECT 3.752 17.569 3.808 17.769 ;
 RECT 4.508 17.4985 4.564 17.6985 ;
 RECT 2.24 17.299 2.296 17.499 ;
 RECT 0.392 18.559 0.448 18.759 ;
 RECT 0.812 18.645 0.868 18.845 ;
 RECT 0.644 18.559 0.7 18.759 ;
 RECT 1.232 18.559 1.288 18.759 ;
 RECT 1.4 18.559 1.456 18.759 ;
 RECT 1.568 18.559 1.624 18.759 ;
 RECT 1.82 18.559 1.876 18.759 ;
 RECT 2.24 18.559 2.296 18.759 ;
 RECT 2.744 18.469 2.8 18.669 ;
 RECT 3.164 18.559 3.22 18.759 ;
 RECT 3.92 18.559 3.976 18.759 ;
 RECT 3.752 18.829 3.808 19.029 ;
 RECT 4.508 18.7585 4.564 18.9585 ;
 RECT 3.5 19.8615 3.556 20.0615 ;
 RECT 0.392 19.819 0.448 20.019 ;
 RECT 0.644 19.819 0.7 20.019 ;
 RECT 1.232 19.819 1.288 20.019 ;
 RECT 0.98 19.7285 1.036 19.9285 ;
 RECT 1.4 19.819 1.456 20.019 ;
 RECT 1.568 19.819 1.624 20.019 ;
 RECT 2.072 19.729 2.128 19.929 ;
 RECT 1.82 19.819 1.876 20.019 ;
 RECT 2.744 19.729 2.8 19.929 ;
 RECT 3.164 19.819 3.22 20.019 ;
 RECT 3.92 19.819 3.976 20.019 ;
 RECT 3.752 20.089 3.808 20.289 ;
 RECT 4.508 20.0185 4.564 20.2185 ;
 RECT 2.24 19.819 2.296 20.019 ;
 END
 END vss.gds1278
 PIN vss.gds1279
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.134 18.1395 10.194 18.3395 ;
 END
 END vss.gds1279
 PIN vss.gds1280
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.966 18.1395 10.026 18.3395 ;
 END
 END vss.gds1280
 PIN vss.gds1281
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.798 18.1395 9.858 18.3395 ;
 END
 END vss.gds1281
 PIN vss.gds1282
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 18.1395 9.69 18.3395 ;
 END
 END vss.gds1282
 PIN vss.gds1283
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.462 18.1395 9.522 18.3395 ;
 END
 END vss.gds1283
 PIN vss.gds1284
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 18.1395 9.018 18.3395 ;
 END
 END vss.gds1284
 PIN vss.gds1285
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.79 18.1395 8.85 18.3395 ;
 END
 END vss.gds1285
 PIN vss.gds1286
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.622 18.1395 8.682 18.3395 ;
 END
 END vss.gds1286
 PIN vss.gds1287
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.454 18.1395 8.514 18.3395 ;
 END
 END vss.gds1287
 PIN vss.gds1288
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 18.5015 5.474 18.7015 ;
 END
 END vss.gds1288
 PIN vss.gds1289
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 18.1395 8.346 18.3395 ;
 END
 END vss.gds1289
 PIN vss.gds1290
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.118 18.1395 8.178 18.3395 ;
 END
 END vss.gds1290
 PIN vss.gds1291
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.95 18.1395 8.01 18.3395 ;
 END
 END vss.gds1291
 PIN vss.gds1292
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.294 18.1395 9.354 18.3395 ;
 END
 END vss.gds1292
 PIN vss.gds1293
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.782 18.1395 7.842 18.3395 ;
 END
 END vss.gds1293
 PIN vss.gds1294
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 18.1395 7.674 18.3395 ;
 END
 END vss.gds1294
 PIN vss.gds1295
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.126 18.1395 9.186 18.3395 ;
 END
 END vss.gds1295
 PIN vss.gds1296
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.446 18.1395 7.506 18.3395 ;
 END
 END vss.gds1296
 PIN vss.gds1297
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.278 18.1395 7.338 18.3395 ;
 END
 END vss.gds1297
 PIN vss.gds1298
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.11 18.1395 7.17 18.3395 ;
 END
 END vss.gds1298
 PIN vss.gds1299
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 18.5015 5.73 18.7015 ;
 END
 END vss.gds1299
 PIN vss.gds1300
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 17.923 5.986 18.123 ;
 END
 END vss.gds1300
 PIN vss.gds1301
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 17.719 6.434 17.919 ;
 END
 END vss.gds1301
 PIN vss.gds1302
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 17.72 6.178 17.92 ;
 END
 END vss.gds1302
 PIN vss.gds1303
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 6.692 17.442 6.748 17.642 ;
 RECT 6.692 16.182 6.748 16.382 ;
 RECT 6.524 16.032 6.58 16.232 ;
 RECT 6.608 16.309 6.664 16.509 ;
 RECT 6.608 17.569 6.664 17.769 ;
 RECT 6.524 17.292 6.58 17.492 ;
 RECT 6.608 18.829 6.664 19.029 ;
 RECT 6.524 18.552 6.58 18.752 ;
 RECT 6.692 18.702 6.748 18.902 ;
 RECT 6.692 19.962 6.748 20.162 ;
 RECT 6.608 20.089 6.664 20.289 ;
 RECT 6.524 19.812 6.58 20.012 ;
 END
 END vss.gds1303
 PIN vss.gds1304
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 20.318 13.898 20.518 ;
 END
 END vss.gds1304
 PIN vss.gds1305
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 16.538 13.898 16.738 ;
 END
 END vss.gds1305
 PIN vss.gds1306
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 16.578 14.87 16.778 ;
 END
 END vss.gds1306
 PIN vss.gds1307
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 19.058 13.898 19.258 ;
 END
 END vss.gds1307
 PIN vss.gds1308
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 19.098 14.87 19.298 ;
 END
 END vss.gds1308
 PIN vss.gds1309
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 17.798 13.898 17.998 ;
 END
 END vss.gds1309
 PIN vss.gds1310
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 17.838 14.87 18.038 ;
 END
 END vss.gds1310
 PIN vss.gds1311
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.15 18.1395 12.21 18.3395 ;
 END
 END vss.gds1311
 PIN vss.gds1312
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.982 18.1395 12.042 18.3395 ;
 END
 END vss.gds1312
 PIN vss.gds1313
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.814 18.1395 11.874 18.3395 ;
 END
 END vss.gds1313
 PIN vss.gds1314
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.478 18.1395 11.538 18.3395 ;
 END
 END vss.gds1314
 PIN vss.gds1315
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.31 18.1395 11.37 18.3395 ;
 END
 END vss.gds1315
 PIN vss.gds1316
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 18.4865 13.058 18.6865 ;
 END
 END vss.gds1316
 PIN vss.gds1317
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 18.1395 11.706 18.3395 ;
 END
 END vss.gds1317
 PIN vss.gds1318
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.142 18.1395 11.202 18.3395 ;
 END
 END vss.gds1318
 PIN vss.gds1319
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.806 18.1395 10.866 18.3395 ;
 END
 END vss.gds1319
 PIN vss.gds1320
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.638 18.1395 10.698 18.3395 ;
 END
 END vss.gds1320
 PIN vss.gds1321
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.47 18.1395 10.53 18.3395 ;
 END
 END vss.gds1321
 PIN vss.gds1322
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 18.1395 11.034 18.3395 ;
 END
 END vss.gds1322
 PIN vss.gds1323
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 18.1395 10.362 18.3395 ;
 END
 END vss.gds1323
 PIN vss.gds1324
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 18.18 15.162 18.38 ;
 END
 END vss.gds1324
 PIN vss.gds1325
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 18.18 14.498 18.38 ;
 END
 END vss.gds1325
 PIN vss.gds1326
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 18.1395 13.658 18.3395 ;
 END
 END vss.gds1326
 PIN vss.gds1327
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.262 18.192 13.318 18.392 ;
 END
 END vss.gds1327
 PIN vss.gds1328
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 18.061 12.378 18.261 ;
 END
 END vss.gds1328
 PIN vss.gds1329
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 18.5015 12.59 18.7015 ;
 END
 END vss.gds1329
 PIN vss.gds1330
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 18.0435 12.818 18.2435 ;
 END
 END vss.gds1330
 PIN vss.gds1331
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 14.336 19.829 14.392 20.029 ;
 RECT 14.168 19.829 14.224 20.029 ;
 RECT 14 19.236 14.056 19.409 ;
 RECT 14.168 19.209 14.224 19.409 ;
 RECT 14 16.716 14.056 16.889 ;
 RECT 14.168 16.689 14.224 16.889 ;
 RECT 14 17.976 14.056 18.149 ;
 RECT 14.168 17.949 14.224 18.149 ;
 RECT 14.336 16.049 14.392 16.249 ;
 RECT 14.168 16.049 14.224 16.249 ;
 RECT 14.336 18.569 14.392 18.769 ;
 RECT 14.168 18.569 14.224 18.769 ;
 RECT 14.336 17.309 14.392 17.509 ;
 RECT 14.168 17.309 14.224 17.509 ;
 RECT 13.664 17.443 13.72 17.643 ;
 RECT 15.008 17.519 15.064 17.719 ;
 RECT 14.84 17.993 14.896 18.158 ;
 RECT 14.672 17.993 14.728 18.158 ;
 RECT 13.664 16.183 13.72 16.383 ;
 RECT 15.008 16.259 15.064 16.459 ;
 RECT 14.84 16.733 14.896 16.898 ;
 RECT 14.672 16.733 14.728 16.898 ;
 RECT 15.008 18.779 15.064 18.979 ;
 RECT 14.84 19.253 14.896 19.418 ;
 RECT 14.672 19.253 14.728 19.418 ;
 RECT 13.664 18.703 13.72 18.903 ;
 RECT 13.664 19.963 13.72 20.163 ;
 RECT 15.008 20.039 15.064 20.239 ;
 RECT 15.176 18.1425 15.232 18.3425 ;
 RECT 12.824 17.9405 12.88 18.1405 ;
 RECT 13.496 18.015 13.552 18.215 ;
 RECT 12.488 17.9775 12.544 18.1775 ;
 RECT 13.328 17.8805 13.384 18.0805 ;
 RECT 13.16 17.9405 13.216 18.1405 ;
 RECT 12.992 17.9405 13.048 18.1405 ;
 RECT 12.656 17.9775 12.712 18.1775 ;
 END
 END vss.gds1331
 PIN vss.gds1332
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 18.553 16.146 18.753 ;
 END
 END vss.gds1332
 PIN vss.gds1333
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 18.036 15.418 18.236 ;
 END
 END vss.gds1333
 PIN vss.gds1334
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 18.1395 20.274 18.3395 ;
 END
 END vss.gds1334
 PIN vss.gds1335
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 19.813 16.146 20.013 ;
 END
 END vss.gds1335
 PIN vss.gds1336
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 18.1395 18.93 18.3395 ;
 END
 END vss.gds1336
 PIN vss.gds1337
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.038 18.1395 19.098 18.3395 ;
 END
 END vss.gds1337
 PIN vss.gds1338
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.206 18.1395 19.266 18.3395 ;
 END
 END vss.gds1338
 PIN vss.gds1339
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.374 18.1395 19.434 18.3395 ;
 END
 END vss.gds1339
 PIN vss.gds1340
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 18.1395 19.602 18.3395 ;
 END
 END vss.gds1340
 PIN vss.gds1341
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 17.293 16.146 17.493 ;
 END
 END vss.gds1341
 PIN vss.gds1342
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 16.033 16.146 16.233 ;
 END
 END vss.gds1342
 PIN vss.gds1343
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 18.0435 17.314 18.2435 ;
 END
 END vss.gds1343
 PIN vss.gds1344
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 18.0985 16.994 18.2985 ;
 END
 END vss.gds1344
 PIN vss.gds1345
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.71 18.1395 19.77 18.3395 ;
 END
 END vss.gds1345
 PIN vss.gds1346
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.878 18.1395 19.938 18.3395 ;
 END
 END vss.gds1346
 PIN vss.gds1347
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 18.18 15.842 18.38 ;
 END
 END vss.gds1347
 PIN vss.gds1348
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 18.192 16.814 18.392 ;
 END
 END vss.gds1348
 PIN vss.gds1349
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.046 18.1395 20.106 18.3395 ;
 END
 END vss.gds1349
 PIN vss.gds1350
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.702 18.1395 18.762 18.3395 ;
 END
 END vss.gds1350
 PIN vss.gds1351
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.534 18.1395 18.594 18.3395 ;
 END
 END vss.gds1351
 PIN vss.gds1352
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.366 18.1395 18.426 18.3395 ;
 END
 END vss.gds1352
 PIN vss.gds1353
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 18.061 18.258 18.261 ;
 END
 END vss.gds1353
 PIN vss.gds1354
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 18.0435 17.834 18.2435 ;
 END
 END vss.gds1354
 PIN vss.gds1355
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.438 18.1955 17.494 18.3955 ;
 END
 END vss.gds1355
 PIN vss.gds1356
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 17.9465 16.49 18.1465 ;
 END
 END vss.gds1356
 PIN vss.gds1357
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.986 17.923 18.026 18.123 ;
 END
 END vss.gds1357
 PIN vss.gds1358
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 15.596 19.48 15.652 19.68 ;
 RECT 15.848 19.483 15.904 19.683 ;
 RECT 15.596 18.22 15.652 18.42 ;
 RECT 15.848 18.223 15.904 18.423 ;
 RECT 16.52 19.256 16.576 19.409 ;
 RECT 15.764 19.253 15.82 19.418 ;
 RECT 15.596 19.253 15.652 19.418 ;
 RECT 15.596 15.7 15.652 15.9 ;
 RECT 15.848 15.703 15.904 15.903 ;
 RECT 16.52 16.736 16.576 16.889 ;
 RECT 15.764 16.733 15.82 16.898 ;
 RECT 15.596 16.733 15.652 16.898 ;
 RECT 15.596 16.96 15.652 17.16 ;
 RECT 15.848 16.963 15.904 17.163 ;
 RECT 16.52 17.996 16.576 18.149 ;
 RECT 15.764 17.993 15.82 18.158 ;
 RECT 15.596 17.993 15.652 18.158 ;
 RECT 16.856 17.3675 16.912 17.5675 ;
 RECT 16.352 17.6195 16.408 17.8195 ;
 RECT 16.352 16.3595 16.408 16.5595 ;
 RECT 16.856 16.1075 16.912 16.3075 ;
 RECT 15.428 17.519 15.484 17.719 ;
 RECT 15.428 16.259 15.484 16.459 ;
 RECT 15.428 18.779 15.484 18.979 ;
 RECT 16.352 18.8795 16.408 19.0795 ;
 RECT 16.856 18.6275 16.912 18.8275 ;
 RECT 15.428 20.039 15.484 20.239 ;
 RECT 16.856 19.8875 16.912 20.0875 ;
 RECT 16.352 20.1395 16.408 20.3395 ;
 RECT 17.864 17.9775 17.92 18.1775 ;
 RECT 17.696 17.979 17.752 18.179 ;
 RECT 17.528 17.9775 17.584 18.1775 ;
 RECT 17.36 17.9775 17.416 18.1775 ;
 RECT 17.192 17.9775 17.248 18.1775 ;
 RECT 18.032 17.9775 18.088 18.1775 ;
 RECT 17.024 18.0915 17.08 18.2915 ;
 END
 END vss.gds1358
 PIN vss.gds1359
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.17 18.1395 25.23 18.3395 ;
 END
 END vss.gds1359
 PIN vss.gds1360
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.002 18.1395 25.062 18.3395 ;
 END
 END vss.gds1360
 PIN vss.gds1361
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.834 18.1395 24.894 18.3395 ;
 END
 END vss.gds1361
 PIN vss.gds1362
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.498 18.1395 24.558 18.3395 ;
 END
 END vss.gds1362
 PIN vss.gds1363
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.33 18.1395 24.39 18.3395 ;
 END
 END vss.gds1363
 PIN vss.gds1364
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.162 18.1395 24.222 18.3395 ;
 END
 END vss.gds1364
 PIN vss.gds1365
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.382 18.1395 20.442 18.3395 ;
 END
 END vss.gds1365
 PIN vss.gds1366
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.55 18.1395 20.61 18.3395 ;
 END
 END vss.gds1366
 PIN vss.gds1367
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.718 18.1395 20.778 18.3395 ;
 END
 END vss.gds1367
 PIN vss.gds1368
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.054 18.1395 21.114 18.3395 ;
 END
 END vss.gds1368
 PIN vss.gds1369
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.222 18.1395 21.282 18.3395 ;
 END
 END vss.gds1369
 PIN vss.gds1370
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.39 18.1395 21.45 18.3395 ;
 END
 END vss.gds1370
 PIN vss.gds1371
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.726 18.1395 21.786 18.3395 ;
 END
 END vss.gds1371
 PIN vss.gds1372
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.894 18.1395 21.954 18.3395 ;
 END
 END vss.gds1372
 PIN vss.gds1373
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.062 18.1395 22.122 18.3395 ;
 END
 END vss.gds1373
 PIN vss.gds1374
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.398 18.1395 22.458 18.3395 ;
 END
 END vss.gds1374
 PIN vss.gds1375
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.566 18.1395 22.626 18.3395 ;
 END
 END vss.gds1375
 PIN vss.gds1376
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.734 18.1395 22.794 18.3395 ;
 END
 END vss.gds1376
 PIN vss.gds1377
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 18.1395 24.726 18.3395 ;
 END
 END vss.gds1377
 PIN vss.gds1378
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 18.1395 21.618 18.3395 ;
 END
 END vss.gds1378
 PIN vss.gds1379
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 18.1395 20.946 18.3395 ;
 END
 END vss.gds1379
 PIN vss.gds1380
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 18.1395 22.29 18.3395 ;
 END
 END vss.gds1380
 PIN vss.gds1381
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 18.1395 22.962 18.3395 ;
 END
 END vss.gds1381
 PIN vss.gds1382
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.07 18.1395 23.13 18.3395 ;
 END
 END vss.gds1382
 PIN vss.gds1383
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.238 18.1395 23.298 18.3395 ;
 END
 END vss.gds1383
 PIN vss.gds1384
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.406 18.1395 23.466 18.3395 ;
 END
 END vss.gds1384
 PIN vss.gds1385
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 18.1395 23.634 18.3395 ;
 END
 END vss.gds1385
 PIN vss.gds1386
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 23.912 17.456 23.968 17.656 ;
 RECT 23.912 16.196 23.968 16.396 ;
 RECT 23.912 18.716 23.968 18.916 ;
 RECT 23.912 19.976 23.968 20.176 ;
 RECT 23.744 18.086 23.8 18.286 ;
 END
 END vss.gds1386
 PIN vss.gds1387
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.202 18.1395 29.262 18.3395 ;
 END
 END vss.gds1387
 PIN vss.gds1388
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.034 18.1395 29.094 18.3395 ;
 END
 END vss.gds1388
 PIN vss.gds1389
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.866 18.1395 28.926 18.3395 ;
 END
 END vss.gds1389
 PIN vss.gds1390
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.53 18.1395 28.59 18.3395 ;
 END
 END vss.gds1390
 PIN vss.gds1391
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.362 18.1395 28.422 18.3395 ;
 END
 END vss.gds1391
 PIN vss.gds1392
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.194 18.1395 28.254 18.3395 ;
 END
 END vss.gds1392
 PIN vss.gds1393
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.858 18.1395 27.918 18.3395 ;
 END
 END vss.gds1393
 PIN vss.gds1394
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.69 18.1395 27.75 18.3395 ;
 END
 END vss.gds1394
 PIN vss.gds1395
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.522 18.1395 27.582 18.3395 ;
 END
 END vss.gds1395
 PIN vss.gds1396
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.186 18.1395 27.246 18.3395 ;
 END
 END vss.gds1396
 PIN vss.gds1397
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.018 18.1395 27.078 18.3395 ;
 END
 END vss.gds1397
 PIN vss.gds1398
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.85 18.1395 26.91 18.3395 ;
 END
 END vss.gds1398
 PIN vss.gds1399
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.514 18.1395 26.574 18.3395 ;
 END
 END vss.gds1399
 PIN vss.gds1400
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.346 18.1395 26.406 18.3395 ;
 END
 END vss.gds1400
 PIN vss.gds1401
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.178 18.1395 26.238 18.3395 ;
 END
 END vss.gds1401
 PIN vss.gds1402
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.842 18.1395 25.902 18.3395 ;
 END
 END vss.gds1402
 PIN vss.gds1403
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.674 18.1395 25.734 18.3395 ;
 END
 END vss.gds1403
 PIN vss.gds1404
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.506 18.1395 25.566 18.3395 ;
 END
 END vss.gds1404
 PIN vss.gds1405
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 18.1395 28.758 18.3395 ;
 END
 END vss.gds1405
 PIN vss.gds1406
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 18.1395 28.086 18.3395 ;
 END
 END vss.gds1406
 PIN vss.gds1407
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 18.1395 27.414 18.3395 ;
 END
 END vss.gds1407
 PIN vss.gds1408
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 18.1395 26.742 18.3395 ;
 END
 END vss.gds1408
 PIN vss.gds1409
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 18.1395 26.07 18.3395 ;
 END
 END vss.gds1409
 PIN vss.gds1410
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 18.1395 25.398 18.3395 ;
 END
 END vss.gds1410
 PIN vss.gds1411
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 18.061 29.43 18.261 ;
 END
 END vss.gds1411
 PIN vss.gds1412
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 18.4865 30.11 18.6865 ;
 END
 END vss.gds1412
 PIN vss.gds1413
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 18.0435 29.87 18.2435 ;
 END
 END vss.gds1413
 PIN vss.gds1414
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 18.5015 29.642 18.7015 ;
 END
 END vss.gds1414
 PIN vss.gds1415
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.876 17.9405 29.932 18.1405 ;
 RECT 30.212 17.9405 30.268 18.1405 ;
 RECT 29.54 17.9775 29.596 18.1775 ;
 RECT 30.044 17.9405 30.1 18.1405 ;
 RECT 29.708 17.9775 29.764 18.1775 ;
 END
 END vss.gds1415
 PIN vss.gds1416
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 20.318 30.95 20.518 ;
 END
 END vss.gds1416
 PIN vss.gds1417
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 16.578 31.922 16.778 ;
 END
 END vss.gds1417
 PIN vss.gds1418
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 19.098 31.922 19.298 ;
 END
 END vss.gds1418
 PIN vss.gds1419
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 17.838 31.922 18.038 ;
 END
 END vss.gds1419
 PIN vss.gds1420
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 16.538 30.95 16.738 ;
 END
 END vss.gds1420
 PIN vss.gds1421
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 17.798 30.95 17.998 ;
 END
 END vss.gds1421
 PIN vss.gds1422
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 19.058 30.95 19.258 ;
 END
 END vss.gds1422
 PIN vss.gds1423
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.314 18.192 30.37 18.392 ;
 END
 END vss.gds1423
 PIN vss.gds1424
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 18.18 32.214 18.38 ;
 END
 END vss.gds1424
 PIN vss.gds1425
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 18.0985 34.046 18.2985 ;
 END
 END vss.gds1425
 PIN vss.gds1426
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 18.1395 30.71 18.3395 ;
 END
 END vss.gds1426
 PIN vss.gds1427
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 19.813 33.198 20.013 ;
 END
 END vss.gds1427
 PIN vss.gds1428
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 18.553 33.198 18.753 ;
 END
 END vss.gds1428
 PIN vss.gds1429
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 17.293 33.198 17.493 ;
 END
 END vss.gds1429
 PIN vss.gds1430
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 16.033 33.198 16.233 ;
 END
 END vss.gds1430
 PIN vss.gds1431
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 18.18 32.894 18.38 ;
 END
 END vss.gds1431
 PIN vss.gds1432
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 17.9465 33.542 18.1465 ;
 END
 END vss.gds1432
 PIN vss.gds1433
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 18.18 31.55 18.38 ;
 END
 END vss.gds1433
 PIN vss.gds1434
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 18.192 33.866 18.392 ;
 END
 END vss.gds1434
 PIN vss.gds1435
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 18.0435 34.886 18.2435 ;
 END
 END vss.gds1435
 PIN vss.gds1436
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.49 18.1955 34.546 18.3955 ;
 END
 END vss.gds1436
 PIN vss.gds1437
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 18.036 32.47 18.236 ;
 END
 END vss.gds1437
 PIN vss.gds1438
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 18.0435 34.366 18.2435 ;
 END
 END vss.gds1438
 PIN vss.gds1439
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.038 17.923 35.078 18.123 ;
 END
 END vss.gds1439
 PIN vss.gds1440
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 32.648 19.48 32.704 19.68 ;
 RECT 32.9 19.483 32.956 19.683 ;
 RECT 31.388 19.829 31.444 20.029 ;
 RECT 31.22 19.829 31.276 20.029 ;
 RECT 30.716 19.963 30.772 20.163 ;
 RECT 32.648 18.22 32.704 18.42 ;
 RECT 32.9 18.223 32.956 18.423 ;
 RECT 33.572 19.256 33.628 19.409 ;
 RECT 31.052 19.236 31.108 19.409 ;
 RECT 31.22 19.209 31.276 19.409 ;
 RECT 32.816 19.253 32.872 19.418 ;
 RECT 32.648 19.253 32.704 19.418 ;
 RECT 31.892 19.253 31.948 19.418 ;
 RECT 31.724 19.253 31.78 19.418 ;
 RECT 33.572 16.736 33.628 16.889 ;
 RECT 31.052 16.716 31.108 16.889 ;
 RECT 31.22 16.689 31.276 16.889 ;
 RECT 32.816 16.733 32.872 16.898 ;
 RECT 32.648 16.733 32.704 16.898 ;
 RECT 31.892 16.733 31.948 16.898 ;
 RECT 31.724 16.733 31.78 16.898 ;
 RECT 33.572 17.996 33.628 18.149 ;
 RECT 31.052 17.976 31.108 18.149 ;
 RECT 31.22 17.949 31.276 18.149 ;
 RECT 32.816 17.993 32.872 18.158 ;
 RECT 32.648 17.993 32.704 18.158 ;
 RECT 31.892 17.993 31.948 18.158 ;
 RECT 31.724 17.993 31.78 18.158 ;
 RECT 32.648 15.7 32.704 15.9 ;
 RECT 32.9 15.703 32.956 15.903 ;
 RECT 32.648 16.96 32.704 17.16 ;
 RECT 32.9 16.963 32.956 17.163 ;
 RECT 31.388 18.569 31.444 18.769 ;
 RECT 31.22 18.569 31.276 18.769 ;
 RECT 32.06 20.039 32.116 20.239 ;
 RECT 32.48 20.039 32.536 20.239 ;
 RECT 32.06 18.779 32.116 18.979 ;
 RECT 30.716 18.703 30.772 18.903 ;
 RECT 32.48 18.779 32.536 18.979 ;
 RECT 31.388 17.309 31.444 17.509 ;
 RECT 31.22 17.309 31.276 17.509 ;
 RECT 33.404 17.6195 33.46 17.8195 ;
 RECT 33.908 17.3675 33.964 17.5675 ;
 RECT 33.404 16.3595 33.46 16.5595 ;
 RECT 33.908 16.1075 33.964 16.3075 ;
 RECT 31.388 16.049 31.444 16.249 ;
 RECT 31.22 16.049 31.276 16.249 ;
 RECT 30.716 17.443 30.772 17.643 ;
 RECT 32.06 17.519 32.116 17.719 ;
 RECT 32.48 17.519 32.536 17.719 ;
 RECT 30.716 16.183 30.772 16.383 ;
 RECT 32.06 16.259 32.116 16.459 ;
 RECT 32.48 16.259 32.536 16.459 ;
 RECT 33.404 18.8795 33.46 19.0795 ;
 RECT 33.908 18.6275 33.964 18.8275 ;
 RECT 30.548 18.015 30.604 18.215 ;
 RECT 33.908 19.8875 33.964 20.0875 ;
 RECT 33.404 20.1395 33.46 20.3395 ;
 RECT 30.38 17.8805 30.436 18.0805 ;
 RECT 32.228 18.1425 32.284 18.3425 ;
 RECT 34.916 17.9775 34.972 18.1775 ;
 RECT 34.748 17.979 34.804 18.179 ;
 RECT 34.58 17.9775 34.636 18.1775 ;
 RECT 34.412 17.9775 34.468 18.1775 ;
 RECT 34.244 17.9775 34.3 18.1775 ;
 RECT 35.084 17.9775 35.14 18.1775 ;
 RECT 34.076 18.0915 34.132 18.2915 ;
 END
 END vss.gds1440
 PIN vss.gds1441
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.122 18.1395 40.182 18.3395 ;
 END
 END vss.gds1441
 PIN vss.gds1442
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.754 18.1395 35.814 18.3395 ;
 END
 END vss.gds1442
 PIN vss.gds1443
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.09 18.1395 36.15 18.3395 ;
 END
 END vss.gds1443
 PIN vss.gds1444
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.258 18.1395 36.318 18.3395 ;
 END
 END vss.gds1444
 PIN vss.gds1445
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.426 18.1395 36.486 18.3395 ;
 END
 END vss.gds1445
 PIN vss.gds1446
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.762 18.1395 36.822 18.3395 ;
 END
 END vss.gds1446
 PIN vss.gds1447
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.93 18.1395 36.99 18.3395 ;
 END
 END vss.gds1447
 PIN vss.gds1448
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.098 18.1395 37.158 18.3395 ;
 END
 END vss.gds1448
 PIN vss.gds1449
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.434 18.1395 37.494 18.3395 ;
 END
 END vss.gds1449
 PIN vss.gds1450
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.602 18.1395 37.662 18.3395 ;
 END
 END vss.gds1450
 PIN vss.gds1451
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.77 18.1395 37.83 18.3395 ;
 END
 END vss.gds1451
 PIN vss.gds1452
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.106 18.1395 38.166 18.3395 ;
 END
 END vss.gds1452
 PIN vss.gds1453
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.274 18.1395 38.334 18.3395 ;
 END
 END vss.gds1453
 PIN vss.gds1454
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 18.1395 36.654 18.3395 ;
 END
 END vss.gds1454
 PIN vss.gds1455
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 18.1395 37.326 18.3395 ;
 END
 END vss.gds1455
 PIN vss.gds1456
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 18.1395 37.998 18.3395 ;
 END
 END vss.gds1456
 PIN vss.gds1457
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.442 18.1395 38.502 18.3395 ;
 END
 END vss.gds1457
 PIN vss.gds1458
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 18.1395 38.67 18.3395 ;
 END
 END vss.gds1458
 PIN vss.gds1459
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.778 18.1395 38.838 18.3395 ;
 END
 END vss.gds1459
 PIN vss.gds1460
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 18.1395 35.982 18.3395 ;
 END
 END vss.gds1460
 PIN vss.gds1461
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.946 18.1395 39.006 18.3395 ;
 END
 END vss.gds1461
 PIN vss.gds1462
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.586 18.1395 35.646 18.3395 ;
 END
 END vss.gds1462
 PIN vss.gds1463
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.45 18.1395 39.51 18.3395 ;
 END
 END vss.gds1463
 PIN vss.gds1464
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.618 18.1395 39.678 18.3395 ;
 END
 END vss.gds1464
 PIN vss.gds1465
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.114 18.1395 39.174 18.3395 ;
 END
 END vss.gds1465
 PIN vss.gds1466
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.786 18.1395 39.846 18.3395 ;
 END
 END vss.gds1466
 PIN vss.gds1467
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 18.1395 40.014 18.3395 ;
 END
 END vss.gds1467
 PIN vss.gds1468
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.418 18.1395 35.478 18.3395 ;
 END
 END vss.gds1468
 PIN vss.gds1469
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 18.061 35.31 18.261 ;
 END
 END vss.gds1469
 PIN vss.gds1470
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 18.1395 39.342 18.3395 ;
 END
 END vss.gds1470
 PIN vss.gds1471
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.91 18.1395 44.97 18.3395 ;
 END
 END vss.gds1471
 PIN vss.gds1472
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.742 18.1395 44.802 18.3395 ;
 END
 END vss.gds1472
 PIN vss.gds1473
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.574 18.1395 44.634 18.3395 ;
 END
 END vss.gds1473
 PIN vss.gds1474
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.238 18.1395 44.298 18.3395 ;
 END
 END vss.gds1474
 PIN vss.gds1475
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.07 18.1395 44.13 18.3395 ;
 END
 END vss.gds1475
 PIN vss.gds1476
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.902 18.1395 43.962 18.3395 ;
 END
 END vss.gds1476
 PIN vss.gds1477
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.566 18.1395 43.626 18.3395 ;
 END
 END vss.gds1477
 PIN vss.gds1478
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.398 18.1395 43.458 18.3395 ;
 END
 END vss.gds1478
 PIN vss.gds1479
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.23 18.1395 43.29 18.3395 ;
 END
 END vss.gds1479
 PIN vss.gds1480
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.894 18.1395 42.954 18.3395 ;
 END
 END vss.gds1480
 PIN vss.gds1481
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.726 18.1395 42.786 18.3395 ;
 END
 END vss.gds1481
 PIN vss.gds1482
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.558 18.1395 42.618 18.3395 ;
 END
 END vss.gds1482
 PIN vss.gds1483
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.222 18.1395 42.282 18.3395 ;
 END
 END vss.gds1483
 PIN vss.gds1484
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.054 18.1395 42.114 18.3395 ;
 END
 END vss.gds1484
 PIN vss.gds1485
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.886 18.1395 41.946 18.3395 ;
 END
 END vss.gds1485
 PIN vss.gds1486
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.55 18.1395 41.61 18.3395 ;
 END
 END vss.gds1486
 PIN vss.gds1487
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.382 18.1395 41.442 18.3395 ;
 END
 END vss.gds1487
 PIN vss.gds1488
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.214 18.1395 41.274 18.3395 ;
 END
 END vss.gds1488
 PIN vss.gds1489
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.29 18.1395 40.35 18.3395 ;
 END
 END vss.gds1489
 PIN vss.gds1490
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.458 18.1395 40.518 18.3395 ;
 END
 END vss.gds1490
 PIN vss.gds1491
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 18.1395 45.138 18.3395 ;
 END
 END vss.gds1491
 PIN vss.gds1492
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 18.1395 44.466 18.3395 ;
 END
 END vss.gds1492
 PIN vss.gds1493
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 18.1395 43.794 18.3395 ;
 END
 END vss.gds1493
 PIN vss.gds1494
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 18.1395 43.122 18.3395 ;
 END
 END vss.gds1494
 PIN vss.gds1495
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 18.1395 42.45 18.3395 ;
 END
 END vss.gds1495
 PIN vss.gds1496
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 18.1395 41.778 18.3395 ;
 END
 END vss.gds1496
 PIN vss.gds1497
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 18.1395 40.686 18.3395 ;
 END
 END vss.gds1497
 PIN vss.gds1498
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 40.964 18.716 41.02 18.916 ;
 RECT 40.964 17.456 41.02 17.656 ;
 RECT 40.964 16.196 41.02 16.396 ;
 RECT 40.964 19.976 41.02 20.176 ;
 RECT 40.796 18.086 40.852 18.286 ;
 END
 END vss.gds1498
 PIN vss.gds1499
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 20.318 48.002 20.518 ;
 END
 END vss.gds1499
 PIN vss.gds1500
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 16.578 48.974 16.778 ;
 END
 END vss.gds1500
 PIN vss.gds1501
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 19.098 48.974 19.298 ;
 END
 END vss.gds1501
 PIN vss.gds1502
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 17.838 48.974 18.038 ;
 END
 END vss.gds1502
 PIN vss.gds1503
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 17.293 50.25 17.493 ;
 END
 END vss.gds1503
 PIN vss.gds1504
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 19.058 48.002 19.258 ;
 END
 END vss.gds1504
 PIN vss.gds1505
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.366 18.192 47.422 18.392 ;
 END
 END vss.gds1505
 PIN vss.gds1506
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.254 18.1395 46.314 18.3395 ;
 END
 END vss.gds1506
 PIN vss.gds1507
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.086 18.1395 46.146 18.3395 ;
 END
 END vss.gds1507
 PIN vss.gds1508
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.918 18.1395 45.978 18.3395 ;
 END
 END vss.gds1508
 PIN vss.gds1509
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.582 18.1395 45.642 18.3395 ;
 END
 END vss.gds1509
 PIN vss.gds1510
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.414 18.1395 45.474 18.3395 ;
 END
 END vss.gds1510
 PIN vss.gds1511
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.246 18.1395 45.306 18.3395 ;
 END
 END vss.gds1511
 PIN vss.gds1512
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 18.4865 47.162 18.6865 ;
 END
 END vss.gds1512
 PIN vss.gds1513
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 18.061 46.482 18.261 ;
 END
 END vss.gds1513
 PIN vss.gds1514
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 18.1395 45.81 18.3395 ;
 END
 END vss.gds1514
 PIN vss.gds1515
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 18.553 50.25 18.753 ;
 END
 END vss.gds1515
 PIN vss.gds1516
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 19.813 50.25 20.013 ;
 END
 END vss.gds1516
 PIN vss.gds1517
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 18.0435 46.922 18.2435 ;
 END
 END vss.gds1517
 PIN vss.gds1518
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 18.5015 46.694 18.7015 ;
 END
 END vss.gds1518
 PIN vss.gds1519
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 18.1395 47.762 18.3395 ;
 END
 END vss.gds1519
 PIN vss.gds1520
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 18.18 49.266 18.38 ;
 END
 END vss.gds1520
 PIN vss.gds1521
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 18.18 48.602 18.38 ;
 END
 END vss.gds1521
 PIN vss.gds1522
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 17.798 48.002 17.998 ;
 END
 END vss.gds1522
 PIN vss.gds1523
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 16.033 50.25 16.233 ;
 END
 END vss.gds1523
 PIN vss.gds1524
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 16.538 48.002 16.738 ;
 END
 END vss.gds1524
 PIN vss.gds1525
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 18.18 49.946 18.38 ;
 END
 END vss.gds1525
 PIN vss.gds1526
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 18.036 49.522 18.236 ;
 END
 END vss.gds1526
 PIN vss.gds1527
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 49.7 19.48 49.756 19.68 ;
 RECT 49.952 19.483 50.008 19.683 ;
 RECT 48.44 19.829 48.496 20.029 ;
 RECT 48.272 19.829 48.328 20.029 ;
 RECT 47.768 19.963 47.824 20.163 ;
 RECT 49.7 18.22 49.756 18.42 ;
 RECT 49.952 18.223 50.008 18.423 ;
 RECT 48.104 19.236 48.16 19.409 ;
 RECT 48.272 19.209 48.328 19.409 ;
 RECT 49.868 19.253 49.924 19.418 ;
 RECT 49.7 19.253 49.756 19.418 ;
 RECT 48.944 19.253 49 19.418 ;
 RECT 48.776 19.253 48.832 19.418 ;
 RECT 48.104 16.716 48.16 16.889 ;
 RECT 48.272 16.689 48.328 16.889 ;
 RECT 49.868 16.733 49.924 16.898 ;
 RECT 49.7 16.733 49.756 16.898 ;
 RECT 48.944 16.733 49 16.898 ;
 RECT 48.776 16.733 48.832 16.898 ;
 RECT 48.104 17.976 48.16 18.149 ;
 RECT 48.272 17.949 48.328 18.149 ;
 RECT 49.868 17.993 49.924 18.158 ;
 RECT 49.7 17.993 49.756 18.158 ;
 RECT 48.944 17.993 49 18.158 ;
 RECT 48.776 17.993 48.832 18.158 ;
 RECT 49.7 15.7 49.756 15.9 ;
 RECT 49.952 15.703 50.008 15.903 ;
 RECT 49.7 16.96 49.756 17.16 ;
 RECT 49.952 16.963 50.008 17.163 ;
 RECT 49.112 20.039 49.168 20.239 ;
 RECT 49.532 20.039 49.588 20.239 ;
 RECT 48.44 18.569 48.496 18.769 ;
 RECT 48.272 18.569 48.328 18.769 ;
 RECT 47.768 18.703 47.824 18.903 ;
 RECT 49.112 18.779 49.168 18.979 ;
 RECT 49.532 18.779 49.588 18.979 ;
 RECT 48.44 17.309 48.496 17.509 ;
 RECT 48.272 17.309 48.328 17.509 ;
 RECT 49.112 17.519 49.168 17.719 ;
 RECT 49.532 17.519 49.588 17.719 ;
 RECT 47.768 17.443 47.824 17.643 ;
 RECT 48.44 16.049 48.496 16.249 ;
 RECT 48.272 16.049 48.328 16.249 ;
 RECT 49.112 16.259 49.168 16.459 ;
 RECT 49.532 16.259 49.588 16.459 ;
 RECT 47.768 16.183 47.824 16.383 ;
 RECT 47.6 18.015 47.656 18.215 ;
 RECT 47.432 17.8805 47.488 18.0805 ;
 RECT 47.264 17.9405 47.32 18.1405 ;
 RECT 46.928 17.9405 46.984 18.1405 ;
 RECT 47.096 17.9405 47.152 18.1405 ;
 RECT 49.28 18.1425 49.336 18.3425 ;
 RECT 46.592 17.9775 46.648 18.1775 ;
 RECT 46.76 17.9775 46.816 18.1775 ;
 END
 END vss.gds1527
 PIN vss.gds1528
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.638 18.1395 52.698 18.3395 ;
 END
 END vss.gds1528
 PIN vss.gds1529
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.806 18.1395 52.866 18.3395 ;
 END
 END vss.gds1529
 PIN vss.gds1530
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.142 18.1395 53.202 18.3395 ;
 END
 END vss.gds1530
 PIN vss.gds1531
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.31 18.1395 53.37 18.3395 ;
 END
 END vss.gds1531
 PIN vss.gds1532
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.478 18.1395 53.538 18.3395 ;
 END
 END vss.gds1532
 PIN vss.gds1533
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.814 18.1395 53.874 18.3395 ;
 END
 END vss.gds1533
 PIN vss.gds1534
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.982 18.1395 54.042 18.3395 ;
 END
 END vss.gds1534
 PIN vss.gds1535
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.15 18.1395 54.21 18.3395 ;
 END
 END vss.gds1535
 PIN vss.gds1536
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.486 18.1395 54.546 18.3395 ;
 END
 END vss.gds1536
 PIN vss.gds1537
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.654 18.1395 54.714 18.3395 ;
 END
 END vss.gds1537
 PIN vss.gds1538
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.822 18.1395 54.882 18.3395 ;
 END
 END vss.gds1538
 PIN vss.gds1539
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.158 18.1395 55.218 18.3395 ;
 END
 END vss.gds1539
 PIN vss.gds1540
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 18.1395 55.05 18.3395 ;
 END
 END vss.gds1540
 PIN vss.gds1541
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 18.1395 54.378 18.3395 ;
 END
 END vss.gds1541
 PIN vss.gds1542
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 18.192 50.918 18.392 ;
 END
 END vss.gds1542
 PIN vss.gds1543
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 18.1395 53.706 18.3395 ;
 END
 END vss.gds1543
 PIN vss.gds1544
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 18.0985 51.098 18.2985 ;
 END
 END vss.gds1544
 PIN vss.gds1545
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 18.1395 53.034 18.3395 ;
 END
 END vss.gds1545
 PIN vss.gds1546
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 18.0435 51.938 18.2435 ;
 END
 END vss.gds1546
 PIN vss.gds1547
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.542 18.1955 51.598 18.3955 ;
 END
 END vss.gds1547
 PIN vss.gds1548
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 18.0435 51.418 18.2435 ;
 END
 END vss.gds1548
 PIN vss.gds1549
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 17.9465 50.594 18.1465 ;
 END
 END vss.gds1549
 PIN vss.gds1550
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.09 17.923 52.13 18.123 ;
 END
 END vss.gds1550
 PIN vss.gds1551
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.47 18.1395 52.53 18.3395 ;
 END
 END vss.gds1551
 PIN vss.gds1552
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 18.061 52.362 18.261 ;
 END
 END vss.gds1552
 PIN vss.gds1553
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 50.624 19.256 50.68 19.409 ;
 RECT 50.624 16.736 50.68 16.889 ;
 RECT 50.624 17.996 50.68 18.149 ;
 RECT 50.456 18.8795 50.512 19.0795 ;
 RECT 50.96 18.6275 51.016 18.8275 ;
 RECT 50.96 17.3675 51.016 17.5675 ;
 RECT 50.456 17.6195 50.512 17.8195 ;
 RECT 50.456 16.3595 50.512 16.5595 ;
 RECT 50.96 16.1075 51.016 16.3075 ;
 RECT 50.96 19.8875 51.016 20.0875 ;
 RECT 50.456 20.1395 50.512 20.3395 ;
 RECT 51.968 17.9775 52.024 18.1775 ;
 RECT 51.8 17.979 51.856 18.179 ;
 RECT 51.632 17.9775 51.688 18.1775 ;
 RECT 51.464 17.9775 51.52 18.1775 ;
 RECT 51.296 17.9775 51.352 18.1775 ;
 RECT 52.136 17.9775 52.192 18.1775 ;
 RECT 51.128 18.0915 51.184 18.2915 ;
 END
 END vss.gds1553
 PIN vss.gds1554
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.946 18.1395 60.006 18.3395 ;
 END
 END vss.gds1554
 PIN vss.gds1555
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.778 18.1395 59.838 18.3395 ;
 END
 END vss.gds1555
 PIN vss.gds1556
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.61 18.1395 59.67 18.3395 ;
 END
 END vss.gds1556
 PIN vss.gds1557
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.274 18.1395 59.334 18.3395 ;
 END
 END vss.gds1557
 PIN vss.gds1558
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.106 18.1395 59.166 18.3395 ;
 END
 END vss.gds1558
 PIN vss.gds1559
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.938 18.1395 58.998 18.3395 ;
 END
 END vss.gds1559
 PIN vss.gds1560
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.602 18.1395 58.662 18.3395 ;
 END
 END vss.gds1560
 PIN vss.gds1561
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.434 18.1395 58.494 18.3395 ;
 END
 END vss.gds1561
 PIN vss.gds1562
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.266 18.1395 58.326 18.3395 ;
 END
 END vss.gds1562
 PIN vss.gds1563
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.326 18.1395 55.386 18.3395 ;
 END
 END vss.gds1563
 PIN vss.gds1564
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.494 18.1395 55.554 18.3395 ;
 END
 END vss.gds1564
 PIN vss.gds1565
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 18.1395 60.174 18.3395 ;
 END
 END vss.gds1565
 PIN vss.gds1566
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 18.1395 59.502 18.3395 ;
 END
 END vss.gds1566
 PIN vss.gds1567
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 18.1395 58.83 18.3395 ;
 END
 END vss.gds1567
 PIN vss.gds1568
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 18.1395 55.722 18.3395 ;
 END
 END vss.gds1568
 PIN vss.gds1569
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.83 18.1395 55.89 18.3395 ;
 END
 END vss.gds1569
 PIN vss.gds1570
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.998 18.1395 56.058 18.3395 ;
 END
 END vss.gds1570
 PIN vss.gds1571
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.166 18.1395 56.226 18.3395 ;
 END
 END vss.gds1571
 PIN vss.gds1572
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 18.1395 56.394 18.3395 ;
 END
 END vss.gds1572
 PIN vss.gds1573
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.502 18.1395 56.562 18.3395 ;
 END
 END vss.gds1573
 PIN vss.gds1574
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.67 18.1395 56.73 18.3395 ;
 END
 END vss.gds1574
 PIN vss.gds1575
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.838 18.1395 56.898 18.3395 ;
 END
 END vss.gds1575
 PIN vss.gds1576
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.342 18.1395 57.402 18.3395 ;
 END
 END vss.gds1576
 PIN vss.gds1577
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.51 18.1395 57.57 18.3395 ;
 END
 END vss.gds1577
 PIN vss.gds1578
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 18.1395 57.738 18.3395 ;
 END
 END vss.gds1578
 PIN vss.gds1579
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.174 18.1395 57.234 18.3395 ;
 END
 END vss.gds1579
 PIN vss.gds1580
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 18.1395 57.066 18.3395 ;
 END
 END vss.gds1580
 PIN vss.gds1581
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 58.016 18.716 58.072 18.916 ;
 RECT 58.016 17.456 58.072 17.656 ;
 RECT 58.016 16.196 58.072 16.396 ;
 RECT 58.016 19.976 58.072 20.176 ;
 RECT 57.848 18.086 57.904 18.286 ;
 END
 END vss.gds1581
 PIN vss.gds1582
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 20.318 65.054 20.518 ;
 END
 END vss.gds1582
 PIN vss.gds1583
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 16.538 65.054 16.738 ;
 END
 END vss.gds1583
 PIN vss.gds1584
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 17.798 65.054 17.998 ;
 END
 END vss.gds1584
 PIN vss.gds1585
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 19.058 65.054 19.258 ;
 END
 END vss.gds1585
 PIN vss.gds1586
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 18.4865 64.214 18.6865 ;
 END
 END vss.gds1586
 PIN vss.gds1587
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.418 18.192 64.474 18.392 ;
 END
 END vss.gds1587
 PIN vss.gds1588
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.306 18.1395 63.366 18.3395 ;
 END
 END vss.gds1588
 PIN vss.gds1589
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.138 18.1395 63.198 18.3395 ;
 END
 END vss.gds1589
 PIN vss.gds1590
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.97 18.1395 63.03 18.3395 ;
 END
 END vss.gds1590
 PIN vss.gds1591
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.634 18.1395 62.694 18.3395 ;
 END
 END vss.gds1591
 PIN vss.gds1592
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.466 18.1395 62.526 18.3395 ;
 END
 END vss.gds1592
 PIN vss.gds1593
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.298 18.1395 62.358 18.3395 ;
 END
 END vss.gds1593
 PIN vss.gds1594
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.962 18.1395 62.022 18.3395 ;
 END
 END vss.gds1594
 PIN vss.gds1595
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.794 18.1395 61.854 18.3395 ;
 END
 END vss.gds1595
 PIN vss.gds1596
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.626 18.1395 61.686 18.3395 ;
 END
 END vss.gds1596
 PIN vss.gds1597
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.29 18.1395 61.35 18.3395 ;
 END
 END vss.gds1597
 PIN vss.gds1598
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.122 18.1395 61.182 18.3395 ;
 END
 END vss.gds1598
 PIN vss.gds1599
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.954 18.1395 61.014 18.3395 ;
 END
 END vss.gds1599
 PIN vss.gds1600
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.618 18.1395 60.678 18.3395 ;
 END
 END vss.gds1600
 PIN vss.gds1601
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.45 18.1395 60.51 18.3395 ;
 END
 END vss.gds1601
 PIN vss.gds1602
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.282 18.1395 60.342 18.3395 ;
 END
 END vss.gds1602
 PIN vss.gds1603
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 18.061 63.534 18.261 ;
 END
 END vss.gds1603
 PIN vss.gds1604
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 18.1395 62.862 18.3395 ;
 END
 END vss.gds1604
 PIN vss.gds1605
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 18.1395 62.19 18.3395 ;
 END
 END vss.gds1605
 PIN vss.gds1606
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 18.1395 61.518 18.3395 ;
 END
 END vss.gds1606
 PIN vss.gds1607
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 18.1395 60.846 18.3395 ;
 END
 END vss.gds1607
 PIN vss.gds1608
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 18.0435 63.974 18.2435 ;
 END
 END vss.gds1608
 PIN vss.gds1609
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 18.5015 63.746 18.7015 ;
 END
 END vss.gds1609
 PIN vss.gds1610
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 18.1395 64.814 18.3395 ;
 END
 END vss.gds1610
 PIN vss.gds1611
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 65.156 19.236 65.212 19.409 ;
 RECT 65.156 16.716 65.212 16.889 ;
 RECT 65.156 17.976 65.212 18.149 ;
 RECT 64.82 19.963 64.876 20.163 ;
 RECT 64.82 18.703 64.876 18.903 ;
 RECT 64.82 17.443 64.876 17.643 ;
 RECT 64.82 16.183 64.876 16.383 ;
 RECT 64.652 18.015 64.708 18.215 ;
 RECT 64.484 17.8805 64.54 18.0805 ;
 RECT 64.316 17.9405 64.372 18.1405 ;
 RECT 64.148 17.9405 64.204 18.1405 ;
 RECT 63.98 17.9405 64.036 18.1405 ;
 RECT 63.644 17.9775 63.7 18.1775 ;
 RECT 63.812 17.9775 63.868 18.1775 ;
 END
 END vss.gds1611
 PIN vss.gds1612
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 16.578 66.026 16.778 ;
 END
 END vss.gds1612
 PIN vss.gds1613
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 19.098 66.026 19.298 ;
 END
 END vss.gds1613
 PIN vss.gds1614
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 17.838 66.026 18.038 ;
 END
 END vss.gds1614
 PIN vss.gds1615
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.69 18.1395 69.75 18.3395 ;
 END
 END vss.gds1615
 PIN vss.gds1616
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.858 18.1395 69.918 18.3395 ;
 END
 END vss.gds1616
 PIN vss.gds1617
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.194 18.1395 70.254 18.3395 ;
 END
 END vss.gds1617
 PIN vss.gds1618
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 18.0985 68.15 18.2985 ;
 END
 END vss.gds1618
 PIN vss.gds1619
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 18.18 66.318 18.38 ;
 END
 END vss.gds1619
 PIN vss.gds1620
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 19.813 67.302 20.013 ;
 END
 END vss.gds1620
 PIN vss.gds1621
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 18.1395 70.086 18.3395 ;
 END
 END vss.gds1621
 PIN vss.gds1622
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 18.553 67.302 18.753 ;
 END
 END vss.gds1622
 PIN vss.gds1623
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 18.18 66.998 18.38 ;
 END
 END vss.gds1623
 PIN vss.gds1624
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 17.293 67.302 17.493 ;
 END
 END vss.gds1624
 PIN vss.gds1625
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 16.033 67.302 16.233 ;
 END
 END vss.gds1625
 PIN vss.gds1626
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 18.18 65.654 18.38 ;
 END
 END vss.gds1626
 PIN vss.gds1627
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 17.9465 67.646 18.1465 ;
 END
 END vss.gds1627
 PIN vss.gds1628
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 18.036 66.574 18.236 ;
 END
 END vss.gds1628
 PIN vss.gds1629
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 18.192 67.97 18.392 ;
 END
 END vss.gds1629
 PIN vss.gds1630
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 18.0435 68.99 18.2435 ;
 END
 END vss.gds1630
 PIN vss.gds1631
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.594 18.1955 68.65 18.3955 ;
 END
 END vss.gds1631
 PIN vss.gds1632
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 18.0435 68.47 18.2435 ;
 END
 END vss.gds1632
 PIN vss.gds1633
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.142 17.923 69.182 18.123 ;
 END
 END vss.gds1633
 PIN vss.gds1634
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.522 18.1395 69.582 18.3395 ;
 END
 END vss.gds1634
 PIN vss.gds1635
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 18.061 69.414 18.261 ;
 END
 END vss.gds1635
 PIN vss.gds1636
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 66.752 19.48 66.808 19.68 ;
 RECT 67.004 19.483 67.06 19.683 ;
 RECT 67.676 19.256 67.732 19.409 ;
 RECT 65.324 19.209 65.38 19.409 ;
 RECT 66.92 19.253 66.976 19.418 ;
 RECT 66.752 19.253 66.808 19.418 ;
 RECT 65.996 19.253 66.052 19.418 ;
 RECT 65.828 19.253 65.884 19.418 ;
 RECT 67.676 16.736 67.732 16.889 ;
 RECT 65.324 16.689 65.38 16.889 ;
 RECT 66.92 16.733 66.976 16.898 ;
 RECT 66.752 16.733 66.808 16.898 ;
 RECT 65.996 16.733 66.052 16.898 ;
 RECT 65.828 16.733 65.884 16.898 ;
 RECT 67.676 17.996 67.732 18.149 ;
 RECT 65.324 17.949 65.38 18.149 ;
 RECT 66.92 17.993 66.976 18.158 ;
 RECT 66.752 17.993 66.808 18.158 ;
 RECT 65.996 17.993 66.052 18.158 ;
 RECT 65.828 17.993 65.884 18.158 ;
 RECT 65.492 19.829 65.548 20.029 ;
 RECT 65.324 19.829 65.38 20.029 ;
 RECT 66.752 15.7 66.808 15.9 ;
 RECT 67.004 15.703 67.06 15.903 ;
 RECT 66.752 16.96 66.808 17.16 ;
 RECT 67.004 16.963 67.06 17.163 ;
 RECT 65.492 17.309 65.548 17.509 ;
 RECT 65.324 17.309 65.38 17.509 ;
 RECT 66.752 18.22 66.808 18.42 ;
 RECT 67.004 18.223 67.06 18.423 ;
 RECT 66.164 20.039 66.22 20.239 ;
 RECT 66.584 20.039 66.64 20.239 ;
 RECT 68.012 18.6275 68.068 18.8275 ;
 RECT 67.508 18.8795 67.564 19.0795 ;
 RECT 66.164 18.779 66.22 18.979 ;
 RECT 66.584 18.779 66.64 18.979 ;
 RECT 65.492 18.569 65.548 18.769 ;
 RECT 65.324 18.569 65.38 18.769 ;
 RECT 66.164 17.519 66.22 17.719 ;
 RECT 66.584 17.519 66.64 17.719 ;
 RECT 67.508 17.6195 67.564 17.8195 ;
 RECT 68.012 17.3675 68.068 17.5675 ;
 RECT 68.012 16.1075 68.068 16.3075 ;
 RECT 67.508 16.3595 67.564 16.5595 ;
 RECT 66.164 16.259 66.22 16.459 ;
 RECT 65.492 16.049 65.548 16.249 ;
 RECT 65.324 16.049 65.38 16.249 ;
 RECT 66.584 16.259 66.64 16.459 ;
 RECT 68.012 19.8875 68.068 20.0875 ;
 RECT 67.508 20.1395 67.564 20.3395 ;
 RECT 66.332 18.1425 66.388 18.3425 ;
 RECT 69.02 17.9775 69.076 18.1775 ;
 RECT 68.852 17.979 68.908 18.179 ;
 RECT 68.684 17.9775 68.74 18.1775 ;
 RECT 68.516 17.9775 68.572 18.1775 ;
 RECT 68.348 17.9775 68.404 18.1775 ;
 RECT 69.188 17.9775 69.244 18.1775 ;
 RECT 68.18 18.0915 68.236 18.2915 ;
 END
 END vss.gds1636
 PIN vss.gds1637
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.362 18.1395 70.422 18.3395 ;
 END
 END vss.gds1637
 PIN vss.gds1638
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.53 18.1395 70.59 18.3395 ;
 END
 END vss.gds1638
 PIN vss.gds1639
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.866 18.1395 70.926 18.3395 ;
 END
 END vss.gds1639
 PIN vss.gds1640
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.034 18.1395 71.094 18.3395 ;
 END
 END vss.gds1640
 PIN vss.gds1641
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.202 18.1395 71.262 18.3395 ;
 END
 END vss.gds1641
 PIN vss.gds1642
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.538 18.1395 71.598 18.3395 ;
 END
 END vss.gds1642
 PIN vss.gds1643
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.706 18.1395 71.766 18.3395 ;
 END
 END vss.gds1643
 PIN vss.gds1644
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.874 18.1395 71.934 18.3395 ;
 END
 END vss.gds1644
 PIN vss.gds1645
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.21 18.1395 72.27 18.3395 ;
 END
 END vss.gds1645
 PIN vss.gds1646
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.378 18.1395 72.438 18.3395 ;
 END
 END vss.gds1646
 PIN vss.gds1647
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.546 18.1395 72.606 18.3395 ;
 END
 END vss.gds1647
 PIN vss.gds1648
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.882 18.1395 72.942 18.3395 ;
 END
 END vss.gds1648
 PIN vss.gds1649
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.05 18.1395 73.11 18.3395 ;
 END
 END vss.gds1649
 PIN vss.gds1650
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 18.1395 71.43 18.3395 ;
 END
 END vss.gds1650
 PIN vss.gds1651
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 18.1395 72.102 18.3395 ;
 END
 END vss.gds1651
 PIN vss.gds1652
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 18.1395 72.774 18.3395 ;
 END
 END vss.gds1652
 PIN vss.gds1653
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 18.1395 70.758 18.3395 ;
 END
 END vss.gds1653
 PIN vss.gds1654
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.554 18.1395 73.614 18.3395 ;
 END
 END vss.gds1654
 PIN vss.gds1655
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.722 18.1395 73.782 18.3395 ;
 END
 END vss.gds1655
 PIN vss.gds1656
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 18.1395 73.446 18.3395 ;
 END
 END vss.gds1656
 PIN vss.gds1657
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.218 18.1395 73.278 18.3395 ;
 END
 END vss.gds1657
 PIN vss.gds1658
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.89 18.1395 73.95 18.3395 ;
 END
 END vss.gds1658
 PIN vss.gds1659
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.394 18.1395 74.454 18.3395 ;
 END
 END vss.gds1659
 PIN vss.gds1660
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 18.1395 74.118 18.3395 ;
 END
 END vss.gds1660
 PIN vss.gds1661
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.562 18.1395 74.622 18.3395 ;
 END
 END vss.gds1661
 PIN vss.gds1662
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 18.1395 74.79 18.3395 ;
 END
 END vss.gds1662
 PIN vss.gds1663
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.226 18.1395 74.286 18.3395 ;
 END
 END vss.gds1663
 PIN vss.gds1664
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.746 24.742 2.802 24.942 ;
 END
 END vss.gds1664
 PIN vss.gds1665
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.646 24.2955 1.702 24.4955 ;
 END
 END vss.gds1665
 PIN vss.gds1666
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.282 22.919 4.338 23.119 ;
 END
 END vss.gds1666
 PIN vss.gds1667
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 22.9435 3.142 23.1435 ;
 END
 END vss.gds1667
 PIN vss.gds1668
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 25.428 4.882 25.628 ;
 END
 END vss.gds1668
 PIN vss.gds1669
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.562 25.371 3.602 25.571 ;
 END
 END vss.gds1669
 PIN vss.gds1670
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 22.8415 0.942 23.0415 ;
 END
 END vss.gds1670
 PIN vss.gds1671
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.286 21.821 3.326 22.021 ;
 END
 END vss.gds1671
 PIN vss.gds1672
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 22.8725 4.194 23.0725 ;
 END
 END vss.gds1672
 PIN vss.gds1673
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 22.444 5.074 22.644 ;
 END
 END vss.gds1673
 PIN vss.gds1674
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 23.4125 0.718 23.6125 ;
 END
 END vss.gds1674
 PIN vss.gds1675
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 21.426 4.882 21.626 ;
 END
 END vss.gds1675
 PIN vss.gds1676
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 22.1335 0.602 22.3335 ;
 END
 END vss.gds1676
 PIN vss.gds1677
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 23.8245 2.122 24.0245 ;
 END
 END vss.gds1677
 PIN vss.gds1678
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 23.5625 1.282 23.7625 ;
 END
 END vss.gds1678
 PIN vss.gds1679
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 23.436 1.462 23.636 ;
 END
 END vss.gds1679
 PIN vss.gds1680
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 23.7605 2.302 23.9605 ;
 END
 END vss.gds1680
 PIN vss.gds1681
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 23.5315 4.002 23.7315 ;
 END
 END vss.gds1681
 PIN vss.gds1682
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 23.6595 5.282 23.8595 ;
 END
 END vss.gds1682
 PIN vss.gds1683
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 23.504 0.29 23.704 ;
 END
 END vss.gds1683
 PIN vss.gds1684
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 3.5 24.765 3.556 24.916 ;
 RECT 3.752 24.765 3.808 24.937 ;
 RECT 2.66 24.778 2.716 24.978 ;
 RECT 3.164 24.498 3.22 24.698 ;
 RECT 3.416 24.535 3.472 24.717 ;
 RECT 4.004 24.6325 4.06 24.8325 ;
 RECT 3.836 24.498 3.892 24.698 ;
 RECT 0.56 24.7975 0.616 24.9975 ;
 RECT 1.568 24.759 1.624 24.959 ;
 RECT 0.98 24.759 1.036 24.959 ;
 RECT 3.164 22.09 3.22 22.29 ;
 RECT 3.416 22.071 3.472 22.253 ;
 RECT 4.004 22.09 4.06 22.29 ;
 RECT 3.836 22.09 3.892 22.29 ;
 RECT 0.56 22.071 0.616 22.271 ;
 RECT 1.568 22.071 1.624 22.271 ;
 RECT 0.98 22.071 1.036 22.271 ;
 RECT 3.164 23.154 3.22 23.354 ;
 RECT 4.508 23.216 4.564 23.367 ;
 RECT 4.76 23.191 4.816 23.373 ;
 RECT 5.18 23.191 5.236 23.373 ;
 RECT 2.24 23.154 2.296 23.354 ;
 RECT 3.164 23.434 3.22 23.634 ;
 RECT 3.416 23.2925 3.472 23.4925 ;
 RECT 4.004 23.294 4.06 23.494 ;
 RECT 3.836 23.294 3.892 23.494 ;
 RECT 4.76 20.727 4.816 20.909 ;
 RECT 4.424 20.748 4.48 20.948 ;
 RECT 5.18 20.727 5.236 20.909 ;
 RECT 4.004 20.748 4.06 20.948 ;
 RECT 3.836 20.727 3.892 20.909 ;
 RECT 3.584 20.748 3.64 20.948 ;
 RECT 3.416 20.748 3.472 20.948 ;
 RECT 0.56 20.727 0.616 20.927 ;
 RECT 1.568 20.727 1.624 20.927 ;
 RECT 0.98 20.727 1.036 20.927 ;
 RECT 1.904 20.748 1.96 20.948 ;
 RECT 2.156 20.748 2.212 20.948 ;
 RECT 2.408 20.748 2.464 20.948 ;
 RECT 2.912 20.748 2.968 20.948 ;
 RECT 2.66 20.748 2.716 20.948 ;
 RECT 3.164 20.748 3.22 20.948 ;
 RECT 0.56 23.4535 0.616 23.6535 ;
 RECT 1.568 23.4535 1.624 23.6535 ;
 RECT 0.98 23.4535 1.036 23.6535 ;
 RECT 2.576 23.415 2.632 23.615 ;
 RECT 0.56 23.173 0.616 23.373 ;
 RECT 1.568 23.173 1.624 23.373 ;
 RECT 0.98 23.173 1.036 23.373 ;
 RECT 2.156 23.3405 2.212 23.5405 ;
 RECT 2.912 23.415 2.968 23.615 ;
 RECT 2.744 23.294 2.8 23.494 ;
 RECT 4.256 23.2925 4.312 23.4925 ;
 RECT 4.676 23.434 4.732 23.634 ;
 RECT 4.424 23.423 4.48 23.623 ;
 RECT 3.584 21.81 3.64 22.01 ;
 RECT 4.004 21.81 4.06 22.01 ;
 RECT 4.256 21.9445 4.312 22.1445 ;
 RECT 4.76 21.9485 4.816 22.1485 ;
 RECT 4.508 21.9445 4.564 22.1445 ;
 RECT 5.18 21.9485 5.236 22.1485 ;
 RECT 0.56 21.829 0.616 22.029 ;
 RECT 1.568 21.829 1.624 22.029 ;
 RECT 0.98 21.829 1.036 22.029 ;
 RECT 3.164 21.81 3.22 22.01 ;
 RECT 2.66 21.95 2.716 22.15 ;
 RECT 2.156 21.95 2.212 22.15 ;
 RECT 0.56 24.478 0.616 24.678 ;
 RECT 1.568 24.478 1.624 24.678 ;
 RECT 0.98 24.478 1.036 24.678 ;
 RECT 2.156 24.638 2.212 24.838 ;
 RECT 2.492 24.5815 2.548 24.7815 ;
 RECT 2.828 24.762 2.884 24.962 ;
 RECT 3.248 24.765 3.304 24.937 ;
 RECT 2.324 24.5815 2.38 24.7815 ;
 RECT 1.988 24.4275 2.044 24.6275 ;
 RECT 1.82 24.478 1.876 24.678 ;
 RECT 4.256 24.6365 4.312 24.8365 ;
 RECT 4.676 24.638 4.732 24.838 ;
 RECT 4.424 24.6325 4.48 24.8325 ;
 END
 END vss.gds1684
 PIN vss.gds1685
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.982 22.185 10.022 22.385 ;
 END
 END vss.gds1685
 PIN vss.gds1686
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.31 22.185 9.35 22.385 ;
 END
 END vss.gds1686
 PIN vss.gds1687
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.638 22.185 8.678 22.385 ;
 END
 END vss.gds1687
 PIN vss.gds1688
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.966 22.185 8.006 22.385 ;
 END
 END vss.gds1688
 PIN vss.gds1689
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.294 22.185 7.334 22.385 ;
 END
 END vss.gds1689
 PIN vss.gds1690
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.778 22.49 9.824 22.69 ;
 END
 END vss.gds1690
 PIN vss.gds1691
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.174 22.6675 10.214 22.8675 ;
 END
 END vss.gds1691
 PIN vss.gds1692
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.106 22.49 9.152 22.69 ;
 END
 END vss.gds1692
 PIN vss.gds1693
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.502 22.6675 9.542 22.8675 ;
 END
 END vss.gds1693
 PIN vss.gds1694
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.434 22.49 8.48 22.69 ;
 END
 END vss.gds1694
 PIN vss.gds1695
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.762 22.49 7.808 22.69 ;
 END
 END vss.gds1695
 PIN vss.gds1696
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.09 22.49 7.136 22.69 ;
 END
 END vss.gds1696
 PIN vss.gds1697
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.83 22.6675 8.87 22.8675 ;
 END
 END vss.gds1697
 PIN vss.gds1698
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.158 22.6675 8.198 22.8675 ;
 END
 END vss.gds1698
 PIN vss.gds1699
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.486 22.6675 7.526 22.8675 ;
 END
 END vss.gds1699
 PIN vss.gds1700
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 23.1945 9.69 23.3945 ;
 END
 END vss.gds1700
 PIN vss.gds1701
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 23.1945 9.018 23.3945 ;
 END
 END vss.gds1701
 PIN vss.gds1702
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.942 23.1945 7.002 23.3945 ;
 END
 END vss.gds1702
 PIN vss.gds1703
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.734 23.8755 6.774 24.0755 ;
 END
 END vss.gds1703
 PIN vss.gds1704
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.606 23.7515 6.646 23.9515 ;
 END
 END vss.gds1704
 PIN vss.gds1705
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 23.296 5.474 23.496 ;
 END
 END vss.gds1705
 PIN vss.gds1706
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 23.1945 8.346 23.3945 ;
 END
 END vss.gds1706
 PIN vss.gds1707
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 23.1945 7.674 23.3945 ;
 END
 END vss.gds1707
 PIN vss.gds1708
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 23.7535 5.73 23.9535 ;
 END
 END vss.gds1708
 PIN vss.gds1709
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 24.0515 5.986 24.2515 ;
 END
 END vss.gds1709
 PIN vss.gds1710
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 23.111 6.434 23.311 ;
 END
 END vss.gds1710
 PIN vss.gds1711
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 21.39 6.178 21.59 ;
 END
 END vss.gds1711
 PIN vss.gds1712
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 6.104 23.154 6.16 23.354 ;
 RECT 5.852 23.154 5.908 23.354 ;
 RECT 5.684 23.154 5.74 23.354 ;
 RECT 6.272 20.748 6.328 20.948 ;
 RECT 6.104 20.748 6.16 20.948 ;
 RECT 5.852 20.748 5.908 20.948 ;
 RECT 5.684 20.748 5.74 20.948 ;
 RECT 9.968 21.19 10.024 21.39 ;
 RECT 9.8 21.19 9.856 21.39 ;
 RECT 10.136 21.19 10.192 21.39 ;
 RECT 9.296 21.19 9.352 21.39 ;
 RECT 9.128 21.19 9.184 21.39 ;
 RECT 9.464 21.19 9.52 21.39 ;
 RECT 9.632 21.181 9.688 21.381 ;
 RECT 8.624 21.19 8.68 21.39 ;
 RECT 8.456 21.19 8.512 21.39 ;
 RECT 8.792 21.19 8.848 21.39 ;
 RECT 8.96 21.181 9.016 21.381 ;
 RECT 7.952 21.19 8.008 21.39 ;
 RECT 7.784 21.19 7.84 21.39 ;
 RECT 8.12 21.19 8.176 21.39 ;
 RECT 8.288 21.181 8.344 21.381 ;
 RECT 6.944 21.181 7 21.381 ;
 RECT 9.632 24.5075 9.688 24.7075 ;
 RECT 8.96 24.5075 9.016 24.7075 ;
 RECT 8.288 24.5075 8.344 24.7075 ;
 RECT 6.944 24.302 7 24.502 ;
 RECT 7.616 24.5075 7.672 24.7075 ;
 RECT 9.968 22.7325 10.024 22.9325 ;
 RECT 9.8 22.7325 9.856 22.9325 ;
 RECT 10.136 22.7325 10.192 22.9325 ;
 RECT 9.296 22.7325 9.352 22.9325 ;
 RECT 9.128 22.7325 9.184 22.9325 ;
 RECT 9.632 22.7325 9.688 22.9325 ;
 RECT 9.464 22.7325 9.52 22.9325 ;
 RECT 8.624 22.7325 8.68 22.9325 ;
 RECT 8.456 22.7325 8.512 22.9325 ;
 RECT 8.96 22.7325 9.016 22.9325 ;
 RECT 8.792 22.7325 8.848 22.9325 ;
 RECT 7.952 22.7325 8.008 22.9325 ;
 RECT 7.784 22.7325 7.84 22.9325 ;
 RECT 8.288 22.7325 8.344 22.9325 ;
 RECT 8.12 22.7325 8.176 22.9325 ;
 RECT 7.28 22.7325 7.336 22.9325 ;
 RECT 6.944 22.7325 7 22.9325 ;
 RECT 7.112 22.7325 7.168 22.9325 ;
 RECT 7.616 22.7325 7.672 22.9325 ;
 RECT 7.448 22.7325 7.504 22.9325 ;
 RECT 7.28 21.19 7.336 21.39 ;
 RECT 7.112 21.19 7.168 21.39 ;
 RECT 7.448 21.19 7.504 21.39 ;
 RECT 7.616 21.181 7.672 21.381 ;
 RECT 6.44 20.748 6.496 20.948 ;
 RECT 5.432 23.434 5.488 23.634 ;
 RECT 5.6 23.434 5.656 23.634 ;
 RECT 5.768 23.434 5.824 23.634 ;
 RECT 5.936 23.434 5.992 23.634 ;
 RECT 6.104 23.434 6.16 23.634 ;
 RECT 6.272 23.294 6.328 23.494 ;
 RECT 6.44 23.294 6.496 23.494 ;
 RECT 6.272 21.95 6.328 22.15 ;
 RECT 6.104 21.95 6.16 22.15 ;
 RECT 5.852 21.95 5.908 22.15 ;
 RECT 5.684 21.95 5.74 22.15 ;
 RECT 6.44 21.81 6.496 22.01 ;
 RECT 6.44 22.09 6.496 22.29 ;
 RECT 5.432 24.638 5.488 24.838 ;
 RECT 5.6 24.638 5.656 24.838 ;
 RECT 5.768 24.638 5.824 24.838 ;
 RECT 5.936 24.638 5.992 24.838 ;
 RECT 6.44 24.638 6.496 24.838 ;
 RECT 6.104 24.638 6.16 24.838 ;
 RECT 6.272 24.638 6.328 24.838 ;
 END
 END vss.gds1712
 PIN vss.gds1713
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.998 22.185 12.038 22.385 ;
 END
 END vss.gds1713
 PIN vss.gds1714
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.326 22.185 11.366 22.385 ;
 END
 END vss.gds1714
 PIN vss.gds1715
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.654 22.185 10.694 22.385 ;
 END
 END vss.gds1715
 PIN vss.gds1716
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.262 21.568 14.318 21.768 ;
 END
 END vss.gds1716
 PIN vss.gds1717
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 21.779 14.87 21.979 ;
 END
 END vss.gds1717
 PIN vss.gds1718
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 21.615 13.058 21.815 ;
 END
 END vss.gds1718
 PIN vss.gds1719
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.422 21.6235 13.478 21.8235 ;
 END
 END vss.gds1719
 PIN vss.gds1720
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.794 22.49 11.84 22.69 ;
 END
 END vss.gds1720
 PIN vss.gds1721
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.19 22.6675 12.23 22.8675 ;
 END
 END vss.gds1721
 PIN vss.gds1722
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.122 22.49 11.168 22.69 ;
 END
 END vss.gds1722
 PIN vss.gds1723
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.518 22.6675 11.558 22.8675 ;
 END
 END vss.gds1723
 PIN vss.gds1724
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.45 22.49 10.496 22.69 ;
 END
 END vss.gds1724
 PIN vss.gds1725
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.846 22.6675 10.886 22.8675 ;
 END
 END vss.gds1725
 PIN vss.gds1726
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 23.1945 11.706 23.3945 ;
 END
 END vss.gds1726
 PIN vss.gds1727
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 23.1945 11.034 23.3945 ;
 END
 END vss.gds1727
 PIN vss.gds1728
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 23.1945 10.362 23.3945 ;
 END
 END vss.gds1728
 PIN vss.gds1729
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 23.1285 15.162 23.3285 ;
 END
 END vss.gds1729
 PIN vss.gds1730
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 23.111 14.498 23.311 ;
 END
 END vss.gds1730
 PIN vss.gds1731
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 23.041 13.658 23.241 ;
 END
 END vss.gds1731
 PIN vss.gds1732
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 23.0545 12.378 23.2545 ;
 END
 END vss.gds1732
 PIN vss.gds1733
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 23.3375 12.59 23.5375 ;
 END
 END vss.gds1733
 PIN vss.gds1734
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 23.041 12.818 23.241 ;
 END
 END vss.gds1734
 PIN vss.gds1735
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 12.74 24.778 12.796 24.978 ;
 RECT 14.252 24.759 14.308 24.941 ;
 RECT 15.092 24.819 15.148 25.019 ;
 RECT 14.756 24.778 14.812 24.978 ;
 RECT 14.504 24.759 14.56 24.941 ;
 RECT 12.656 22.09 12.712 22.29 ;
 RECT 13.244 22.071 13.3 22.253 ;
 RECT 12.656 21.81 12.712 22.01 ;
 RECT 13.244 21.847 13.3 22.029 ;
 RECT 13.916 21.95 13.972 22.15 ;
 RECT 13.496 23.154 13.552 23.354 ;
 RECT 13.076 23.154 13.132 23.354 ;
 RECT 13.916 23.154 13.972 23.354 ;
 RECT 14.336 23.154 14.392 23.354 ;
 RECT 14.84 23.154 14.896 23.354 ;
 RECT 14.672 23.191 14.728 23.373 ;
 RECT 15.176 23.0835 15.232 23.2835 ;
 RECT 14.672 23.415 14.728 23.597 ;
 RECT 14.84 23.434 14.896 23.634 ;
 RECT 13.58 20.748 13.636 20.948 ;
 RECT 12.908 20.748 12.964 20.948 ;
 RECT 13.916 20.748 13.972 20.948 ;
 RECT 14.252 20.748 14.308 20.948 ;
 RECT 14.588 20.748 14.644 20.948 ;
 RECT 14.924 20.748 14.98 20.948 ;
 RECT 13.244 20.709 13.3 20.909 ;
 RECT 11.984 21.19 12.04 21.39 ;
 RECT 12.32 21.181 12.376 21.381 ;
 RECT 11.312 21.19 11.368 21.39 ;
 RECT 11.144 21.19 11.2 21.39 ;
 RECT 11.48 21.19 11.536 21.39 ;
 RECT 11.648 21.181 11.704 21.381 ;
 RECT 10.64 21.19 10.696 21.39 ;
 RECT 10.472 21.19 10.528 21.39 ;
 RECT 10.808 21.19 10.864 21.39 ;
 RECT 10.976 21.181 11.032 21.381 ;
 RECT 10.304 21.181 10.36 21.381 ;
 RECT 14 20.496 14.056 20.669 ;
 RECT 14.168 20.469 14.224 20.669 ;
 RECT 13.076 23.5045 13.132 23.7045 ;
 RECT 13.496 23.5045 13.552 23.7045 ;
 RECT 13.916 23.5045 13.972 23.7045 ;
 RECT 14.336 23.5045 14.392 23.7045 ;
 RECT 15.176 23.5045 15.232 23.7045 ;
 RECT 13.244 24.638 13.3 24.838 ;
 RECT 14.252 24.535 14.308 24.717 ;
 RECT 13.916 24.638 13.972 24.838 ;
 RECT 15.092 24.498 15.148 24.698 ;
 RECT 14.756 24.498 14.812 24.698 ;
 RECT 14.588 24.535 14.644 24.717 ;
 RECT 12.32 24.5075 12.376 24.7075 ;
 RECT 11.648 24.5075 11.704 24.7075 ;
 RECT 10.976 24.5075 11.032 24.7075 ;
 RECT 10.304 24.5075 10.36 24.7075 ;
 RECT 11.984 22.7325 12.04 22.9325 ;
 RECT 11.816 22.7325 11.872 22.9325 ;
 RECT 12.32 22.7325 12.376 22.9325 ;
 RECT 12.152 22.7325 12.208 22.9325 ;
 RECT 11.312 22.7325 11.368 22.9325 ;
 RECT 11.144 22.7325 11.2 22.9325 ;
 RECT 11.648 22.7325 11.704 22.9325 ;
 RECT 11.48 22.7325 11.536 22.9325 ;
 RECT 10.64 22.7325 10.696 22.9325 ;
 RECT 10.472 22.7325 10.528 22.9325 ;
 RECT 10.976 22.7325 11.032 22.9325 ;
 RECT 10.808 22.7325 10.864 22.9325 ;
 RECT 10.304 22.7325 10.36 22.9325 ;
 RECT 14.84 20.513 14.896 20.678 ;
 RECT 14.672 20.513 14.728 20.678 ;
 RECT 11.816 21.19 11.872 21.39 ;
 RECT 12.152 21.19 12.208 21.39 ;
 RECT 15.176 20.554 15.232 20.754 ;
 RECT 12.824 20.543 12.88 20.743 ;
 RECT 12.488 20.543 12.544 20.743 ;
 RECT 13.328 20.543 13.384 20.743 ;
 RECT 13.16 20.543 13.216 20.743 ;
 RECT 12.992 20.543 13.048 20.743 ;
 RECT 12.656 20.626 12.712 20.826 ;
 END
 END vss.gds1735
 PIN vss.gds1736
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.894 22.185 19.934 22.385 ;
 END
 END vss.gds1736
 PIN vss.gds1737
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.222 22.185 19.262 22.385 ;
 END
 END vss.gds1737
 PIN vss.gds1738
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.69 22.49 19.736 22.69 ;
 END
 END vss.gds1738
 PIN vss.gds1739
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.086 22.6675 20.126 22.8675 ;
 END
 END vss.gds1739
 PIN vss.gds1740
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 21.568 15.418 21.768 ;
 END
 END vss.gds1740
 PIN vss.gds1741
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 23.1945 20.274 23.3945 ;
 END
 END vss.gds1741
 PIN vss.gds1742
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.17 24.6335 16.226 24.8335 ;
 END
 END vss.gds1742
 PIN vss.gds1743
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.594 25.031 16.65 25.231 ;
 END
 END vss.gds1743
 PIN vss.gds1744
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 24.37 17.314 24.57 ;
 END
 END vss.gds1744
 PIN vss.gds1745
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 23.2245 16.146 23.4245 ;
 END
 END vss.gds1745
 PIN vss.gds1746
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.018 22.49 19.064 22.69 ;
 END
 END vss.gds1746
 PIN vss.gds1747
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.414 22.6675 19.454 22.8675 ;
 END
 END vss.gds1747
 PIN vss.gds1748
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.346 22.49 18.392 22.69 ;
 END
 END vss.gds1748
 PIN vss.gds1749
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.742 22.6675 18.782 22.8675 ;
 END
 END vss.gds1749
 PIN vss.gds1750
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.598 23.595 17.654 23.795 ;
 END
 END vss.gds1750
 PIN vss.gds1751
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.55 22.185 18.59 22.385 ;
 END
 END vss.gds1751
 PIN vss.gds1752
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 23.1945 18.93 23.3945 ;
 END
 END vss.gds1752
 PIN vss.gds1753
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 23.1945 19.602 23.3945 ;
 END
 END vss.gds1753
 PIN vss.gds1754
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 20.957 17.314 21.157 ;
 END
 END vss.gds1754
 PIN vss.gds1755
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 23.2295 16.994 23.4295 ;
 END
 END vss.gds1755
 PIN vss.gds1756
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 23.427 15.842 23.627 ;
 END
 END vss.gds1756
 PIN vss.gds1757
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 21.426 16.814 21.626 ;
 END
 END vss.gds1757
 PIN vss.gds1758
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 23.1945 18.258 23.3945 ;
 END
 END vss.gds1758
 PIN vss.gds1759
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 23.2755 17.834 23.4755 ;
 END
 END vss.gds1759
 PIN vss.gds1760
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 23.128 16.49 23.328 ;
 END
 END vss.gds1760
 PIN vss.gds1761
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 15.428 24.778 15.484 24.978 ;
 RECT 16.016 24.778 16.072 24.978 ;
 RECT 15.848 24.778 15.904 24.978 ;
 RECT 16.52 24.759 16.576 24.941 ;
 RECT 16.268 24.759 16.324 24.941 ;
 RECT 17.108 24.778 17.164 24.978 ;
 RECT 17.276 24.778 17.332 24.978 ;
 RECT 15.932 22.09 15.988 22.29 ;
 RECT 15.764 22.09 15.82 22.29 ;
 RECT 15.596 22.09 15.652 22.29 ;
 RECT 15.428 22.09 15.484 22.29 ;
 RECT 16.604 22.09 16.66 22.29 ;
 RECT 16.184 22.072 16.24 22.249 ;
 RECT 15.932 21.81 15.988 22.01 ;
 RECT 15.764 21.81 15.82 22.01 ;
 RECT 15.596 21.81 15.652 22.01 ;
 RECT 15.428 21.81 15.484 22.01 ;
 RECT 16.184 21.851 16.24 22.029 ;
 RECT 16.352 21.847 16.408 22.047 ;
 RECT 16.688 21.81 16.744 22.01 ;
 RECT 16.1 23.195 16.156 23.367 ;
 RECT 15.848 23.195 15.904 23.367 ;
 RECT 15.512 23.154 15.568 23.354 ;
 RECT 16.52 23.154 16.576 23.354 ;
 RECT 17.528 23.154 17.584 23.354 ;
 RECT 17.024 23.154 17.08 23.354 ;
 RECT 16.1 23.415 16.156 23.593 ;
 RECT 15.512 23.434 15.568 23.634 ;
 RECT 15.848 23.415 15.904 23.593 ;
 RECT 16.604 23.434 16.66 23.634 ;
 RECT 17.108 23.434 17.164 23.634 ;
 RECT 17.528 23.434 17.584 23.634 ;
 RECT 15.932 20.748 15.988 20.948 ;
 RECT 16.268 20.748 16.324 20.948 ;
 RECT 16.604 20.748 16.66 20.948 ;
 RECT 16.94 20.748 16.996 20.948 ;
 RECT 16.52 20.516 16.576 20.669 ;
 RECT 15.764 20.513 15.82 20.678 ;
 RECT 15.596 20.513 15.652 20.678 ;
 RECT 19.88 21.19 19.936 21.39 ;
 RECT 19.712 21.19 19.768 21.39 ;
 RECT 20.048 21.19 20.104 21.39 ;
 RECT 20.216 21.181 20.272 21.381 ;
 RECT 19.208 21.19 19.264 21.39 ;
 RECT 19.04 21.19 19.096 21.39 ;
 RECT 19.376 21.19 19.432 21.39 ;
 RECT 19.544 21.181 19.6 21.381 ;
 RECT 18.2 21.181 18.256 21.381 ;
 RECT 17.276 20.709 17.332 20.909 ;
 RECT 18.536 21.19 18.592 21.39 ;
 RECT 18.368 21.19 18.424 21.39 ;
 RECT 18.704 21.19 18.76 21.39 ;
 RECT 18.872 21.181 18.928 21.381 ;
 RECT 17.78 24.8485 17.836 25.0485 ;
 RECT 16.1 24.535 16.156 24.717 ;
 RECT 15.428 24.498 15.484 24.698 ;
 RECT 15.764 24.535 15.82 24.717 ;
 RECT 16.604 24.498 16.66 24.698 ;
 RECT 17.192 24.535 17.248 24.717 ;
 RECT 20.216 24.5075 20.272 24.7075 ;
 RECT 19.544 24.5075 19.6 24.7075 ;
 RECT 18.2 24.302 18.256 24.502 ;
 RECT 18.872 24.5075 18.928 24.7075 ;
 RECT 19.88 22.7325 19.936 22.9325 ;
 RECT 19.712 22.7325 19.768 22.9325 ;
 RECT 20.216 22.7325 20.272 22.9325 ;
 RECT 20.048 22.7325 20.104 22.9325 ;
 RECT 19.208 22.7325 19.264 22.9325 ;
 RECT 19.04 22.7325 19.096 22.9325 ;
 RECT 19.544 22.7325 19.6 22.9325 ;
 RECT 19.376 22.7325 19.432 22.9325 ;
 RECT 18.536 22.7325 18.592 22.9325 ;
 RECT 18.2 22.7325 18.256 22.9325 ;
 RECT 18.368 22.7325 18.424 22.9325 ;
 RECT 18.872 22.7325 18.928 22.9325 ;
 RECT 18.704 22.7325 18.76 22.9325 ;
 RECT 17.864 20.543 17.92 20.743 ;
 RECT 17.696 20.543 17.752 20.743 ;
 RECT 17.528 20.543 17.584 20.743 ;
 RECT 17.36 20.543 17.416 20.743 ;
 RECT 17.192 20.543 17.248 20.743 ;
 RECT 18.032 20.543 18.088 20.743 ;
 RECT 17.024 20.554 17.08 20.754 ;
 RECT 17.78 22.131 17.836 22.331 ;
 RECT 17.528 22.0615 17.584 22.2615 ;
 RECT 16.94 21.95 16.996 22.15 ;
 RECT 17.276 21.95 17.332 22.15 ;
 RECT 17.108 21.95 17.164 22.15 ;
 RECT 17.864 21.81 17.92 22.01 ;
 END
 END vss.gds1761
 PIN vss.gds1762
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.018 22.185 25.058 22.385 ;
 END
 END vss.gds1762
 PIN vss.gds1763
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.346 22.185 24.386 22.385 ;
 END
 END vss.gds1763
 PIN vss.gds1764
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.254 22.185 23.294 22.385 ;
 END
 END vss.gds1764
 PIN vss.gds1765
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.582 22.185 22.622 22.385 ;
 END
 END vss.gds1765
 PIN vss.gds1766
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.91 22.185 21.95 22.385 ;
 END
 END vss.gds1766
 PIN vss.gds1767
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.238 22.185 21.278 22.385 ;
 END
 END vss.gds1767
 PIN vss.gds1768
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.566 22.185 20.606 22.385 ;
 END
 END vss.gds1768
 PIN vss.gds1769
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.814 22.49 24.86 22.69 ;
 END
 END vss.gds1769
 PIN vss.gds1770
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.21 22.6675 25.25 22.8675 ;
 END
 END vss.gds1770
 PIN vss.gds1771
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.142 22.49 24.188 22.69 ;
 END
 END vss.gds1771
 PIN vss.gds1772
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.538 22.6675 24.578 22.8675 ;
 END
 END vss.gds1772
 PIN vss.gds1773
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.05 22.49 23.096 22.69 ;
 END
 END vss.gds1773
 PIN vss.gds1774
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.446 22.6675 23.486 22.8675 ;
 END
 END vss.gds1774
 PIN vss.gds1775
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.378 22.49 22.424 22.69 ;
 END
 END vss.gds1775
 PIN vss.gds1776
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.774 22.6675 22.814 22.8675 ;
 END
 END vss.gds1776
 PIN vss.gds1777
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.706 22.49 21.752 22.69 ;
 END
 END vss.gds1777
 PIN vss.gds1778
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.102 22.6675 22.142 22.8675 ;
 END
 END vss.gds1778
 PIN vss.gds1779
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.034 22.49 21.08 22.69 ;
 END
 END vss.gds1779
 PIN vss.gds1780
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.43 22.6675 21.47 22.8675 ;
 END
 END vss.gds1780
 PIN vss.gds1781
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.362 22.49 20.408 22.69 ;
 END
 END vss.gds1781
 PIN vss.gds1782
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.758 22.6675 20.798 22.8675 ;
 END
 END vss.gds1782
 PIN vss.gds1783
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.722 23.932 23.762 24.132 ;
 END
 END vss.gds1783
 PIN vss.gds1784
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.866 23.932 23.906 24.132 ;
 END
 END vss.gds1784
 PIN vss.gds1785
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 23.1945 24.726 23.3945 ;
 END
 END vss.gds1785
 PIN vss.gds1786
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 23.1945 21.618 23.3945 ;
 END
 END vss.gds1786
 PIN vss.gds1787
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.994 23.2565 24.054 23.4565 ;
 END
 END vss.gds1787
 PIN vss.gds1788
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 23.1945 20.946 23.3945 ;
 END
 END vss.gds1788
 PIN vss.gds1789
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 23.1945 22.29 23.3945 ;
 END
 END vss.gds1789
 PIN vss.gds1790
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 23.1945 22.962 23.3945 ;
 END
 END vss.gds1790
 PIN vss.gds1791
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 23.2565 23.634 23.4565 ;
 END
 END vss.gds1791
 PIN vss.gds1792
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 25.004 21.19 25.06 21.39 ;
 RECT 24.836 21.19 24.892 21.39 ;
 RECT 25.172 21.19 25.228 21.39 ;
 RECT 24.668 21.181 24.724 21.381 ;
 RECT 23.996 21.0105 24.052 21.2105 ;
 RECT 24.332 21.19 24.388 21.39 ;
 RECT 24.164 21.19 24.22 21.39 ;
 RECT 24.5 21.19 24.556 21.39 ;
 RECT 23.24 21.19 23.296 21.39 ;
 RECT 23.072 21.19 23.128 21.39 ;
 RECT 23.408 21.19 23.464 21.39 ;
 RECT 23.576 21.181 23.632 21.381 ;
 RECT 22.568 21.19 22.624 21.39 ;
 RECT 22.4 21.19 22.456 21.39 ;
 RECT 22.736 21.19 22.792 21.39 ;
 RECT 22.904 21.181 22.96 21.381 ;
 RECT 21.896 21.19 21.952 21.39 ;
 RECT 21.728 21.19 21.784 21.39 ;
 RECT 22.064 21.19 22.12 21.39 ;
 RECT 22.232 21.181 22.288 21.381 ;
 RECT 21.224 21.19 21.28 21.39 ;
 RECT 21.056 21.19 21.112 21.39 ;
 RECT 21.392 21.19 21.448 21.39 ;
 RECT 21.56 21.181 21.616 21.381 ;
 RECT 20.888 21.181 20.944 21.381 ;
 RECT 20.552 21.19 20.608 21.39 ;
 RECT 20.72 21.19 20.776 21.39 ;
 RECT 20.384 21.19 20.44 21.39 ;
 RECT 23.996 24.302 24.052 24.502 ;
 RECT 24.668 24.5075 24.724 24.7075 ;
 RECT 23.576 24.5075 23.632 24.7075 ;
 RECT 22.904 24.5075 22.96 24.7075 ;
 RECT 22.232 24.5075 22.288 24.7075 ;
 RECT 21.56 24.5075 21.616 24.7075 ;
 RECT 20.888 24.5075 20.944 24.7075 ;
 RECT 25.004 22.7325 25.06 22.9325 ;
 RECT 24.836 22.7325 24.892 22.9325 ;
 RECT 25.172 22.7325 25.228 22.9325 ;
 RECT 24.332 22.7325 24.388 22.9325 ;
 RECT 23.996 22.7325 24.052 22.9325 ;
 RECT 24.164 22.7325 24.22 22.9325 ;
 RECT 24.668 22.7325 24.724 22.9325 ;
 RECT 24.5 22.7325 24.556 22.9325 ;
 RECT 23.24 22.7325 23.296 22.9325 ;
 RECT 23.072 22.7325 23.128 22.9325 ;
 RECT 23.576 22.7325 23.632 22.9325 ;
 RECT 23.408 22.7325 23.464 22.9325 ;
 RECT 22.568 22.7325 22.624 22.9325 ;
 RECT 22.4 22.7325 22.456 22.9325 ;
 RECT 22.904 22.7325 22.96 22.9325 ;
 RECT 22.736 22.7325 22.792 22.9325 ;
 RECT 21.896 22.7325 21.952 22.9325 ;
 RECT 21.728 22.7325 21.784 22.9325 ;
 RECT 22.232 22.7325 22.288 22.9325 ;
 RECT 22.064 22.7325 22.12 22.9325 ;
 RECT 21.224 22.7325 21.28 22.9325 ;
 RECT 21.056 22.7325 21.112 22.9325 ;
 RECT 21.56 22.7325 21.616 22.9325 ;
 RECT 21.392 22.7325 21.448 22.9325 ;
 RECT 20.552 22.7325 20.608 22.9325 ;
 RECT 20.888 22.7325 20.944 22.9325 ;
 RECT 20.72 22.7325 20.776 22.9325 ;
 RECT 20.384 22.7325 20.44 22.9325 ;
 RECT 23.744 22.7795 23.8 22.9795 ;
 END
 END vss.gds1792
 PIN vss.gds1793
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.05 22.185 29.09 22.385 ;
 END
 END vss.gds1793
 PIN vss.gds1794
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.378 22.185 28.418 22.385 ;
 END
 END vss.gds1794
 PIN vss.gds1795
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.706 22.185 27.746 22.385 ;
 END
 END vss.gds1795
 PIN vss.gds1796
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.034 22.185 27.074 22.385 ;
 END
 END vss.gds1796
 PIN vss.gds1797
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.362 22.185 26.402 22.385 ;
 END
 END vss.gds1797
 PIN vss.gds1798
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.69 22.185 25.73 22.385 ;
 END
 END vss.gds1798
 PIN vss.gds1799
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.846 22.49 28.892 22.69 ;
 END
 END vss.gds1799
 PIN vss.gds1800
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.242 22.6675 29.282 22.8675 ;
 END
 END vss.gds1800
 PIN vss.gds1801
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.174 22.49 28.22 22.69 ;
 END
 END vss.gds1801
 PIN vss.gds1802
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.57 22.6675 28.61 22.8675 ;
 END
 END vss.gds1802
 PIN vss.gds1803
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.502 22.49 27.548 22.69 ;
 END
 END vss.gds1803
 PIN vss.gds1804
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.898 22.6675 27.938 22.8675 ;
 END
 END vss.gds1804
 PIN vss.gds1805
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.83 22.49 26.876 22.69 ;
 END
 END vss.gds1805
 PIN vss.gds1806
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.226 22.6675 27.266 22.8675 ;
 END
 END vss.gds1806
 PIN vss.gds1807
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.158 22.49 26.204 22.69 ;
 END
 END vss.gds1807
 PIN vss.gds1808
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.554 22.6675 26.594 22.8675 ;
 END
 END vss.gds1808
 PIN vss.gds1809
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.486 22.49 25.532 22.69 ;
 END
 END vss.gds1809
 PIN vss.gds1810
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.882 22.6675 25.922 22.8675 ;
 END
 END vss.gds1810
 PIN vss.gds1811
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 23.1945 28.758 23.3945 ;
 END
 END vss.gds1811
 PIN vss.gds1812
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 23.1945 28.086 23.3945 ;
 END
 END vss.gds1812
 PIN vss.gds1813
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 23.1945 27.414 23.3945 ;
 END
 END vss.gds1813
 PIN vss.gds1814
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 23.1945 26.742 23.3945 ;
 END
 END vss.gds1814
 PIN vss.gds1815
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 23.1945 26.07 23.3945 ;
 END
 END vss.gds1815
 PIN vss.gds1816
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 23.1945 25.398 23.3945 ;
 END
 END vss.gds1816
 PIN vss.gds1817
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 23.0545 29.43 23.2545 ;
 END
 END vss.gds1817
 PIN vss.gds1818
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 21.615 30.11 21.815 ;
 END
 END vss.gds1818
 PIN vss.gds1819
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 23.041 29.87 23.241 ;
 END
 END vss.gds1819
 PIN vss.gds1820
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 23.3375 29.642 23.5375 ;
 END
 END vss.gds1820
 PIN vss.gds1821
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.792 24.778 29.848 24.978 ;
 RECT 29.708 22.09 29.764 22.29 ;
 RECT 29.708 21.81 29.764 22.01 ;
 RECT 30.128 23.154 30.184 23.354 ;
 RECT 29.96 20.748 30.016 20.948 ;
 RECT 30.128 23.5045 30.184 23.7045 ;
 RECT 29.036 21.19 29.092 21.39 ;
 RECT 28.868 21.19 28.924 21.39 ;
 RECT 29.204 21.19 29.26 21.39 ;
 RECT 29.372 21.181 29.428 21.381 ;
 RECT 28.364 21.19 28.42 21.39 ;
 RECT 28.196 21.19 28.252 21.39 ;
 RECT 28.532 21.19 28.588 21.39 ;
 RECT 28.7 21.181 28.756 21.381 ;
 RECT 27.692 21.19 27.748 21.39 ;
 RECT 27.524 21.19 27.58 21.39 ;
 RECT 27.86 21.19 27.916 21.39 ;
 RECT 28.028 21.181 28.084 21.381 ;
 RECT 27.02 21.19 27.076 21.39 ;
 RECT 26.852 21.19 26.908 21.39 ;
 RECT 27.188 21.19 27.244 21.39 ;
 RECT 27.356 21.181 27.412 21.381 ;
 RECT 26.348 21.19 26.404 21.39 ;
 RECT 26.18 21.19 26.236 21.39 ;
 RECT 26.516 21.19 26.572 21.39 ;
 RECT 26.684 21.181 26.74 21.381 ;
 RECT 25.676 21.19 25.732 21.39 ;
 RECT 25.508 21.19 25.564 21.39 ;
 RECT 25.844 21.19 25.9 21.39 ;
 RECT 26.012 21.181 26.068 21.381 ;
 RECT 25.34 21.181 25.396 21.381 ;
 RECT 29.372 24.5075 29.428 24.7075 ;
 RECT 28.7 24.5075 28.756 24.7075 ;
 RECT 28.028 24.5075 28.084 24.7075 ;
 RECT 27.356 24.5075 27.412 24.7075 ;
 RECT 26.684 24.5075 26.74 24.7075 ;
 RECT 26.012 24.5075 26.068 24.7075 ;
 RECT 25.34 24.5075 25.396 24.7075 ;
 RECT 29.036 22.7325 29.092 22.9325 ;
 RECT 28.868 22.7325 28.924 22.9325 ;
 RECT 29.372 22.7325 29.428 22.9325 ;
 RECT 29.204 22.7325 29.26 22.9325 ;
 RECT 28.364 22.7325 28.42 22.9325 ;
 RECT 28.196 22.7325 28.252 22.9325 ;
 RECT 28.7 22.7325 28.756 22.9325 ;
 RECT 28.532 22.7325 28.588 22.9325 ;
 RECT 27.692 22.7325 27.748 22.9325 ;
 RECT 27.524 22.7325 27.58 22.9325 ;
 RECT 28.028 22.7325 28.084 22.9325 ;
 RECT 27.86 22.7325 27.916 22.9325 ;
 RECT 27.02 22.7325 27.076 22.9325 ;
 RECT 26.852 22.7325 26.908 22.9325 ;
 RECT 27.356 22.7325 27.412 22.9325 ;
 RECT 27.188 22.7325 27.244 22.9325 ;
 RECT 26.348 22.7325 26.404 22.9325 ;
 RECT 26.18 22.7325 26.236 22.9325 ;
 RECT 26.684 22.7325 26.74 22.9325 ;
 RECT 26.516 22.7325 26.572 22.9325 ;
 RECT 25.676 22.7325 25.732 22.9325 ;
 RECT 25.508 22.7325 25.564 22.9325 ;
 RECT 26.012 22.7325 26.068 22.9325 ;
 RECT 25.844 22.7325 25.9 22.9325 ;
 RECT 25.34 22.7325 25.396 22.9325 ;
 RECT 29.876 20.543 29.932 20.743 ;
 RECT 30.212 20.543 30.268 20.743 ;
 RECT 29.54 20.543 29.596 20.743 ;
 RECT 30.044 20.543 30.1 20.743 ;
 RECT 29.708 20.626 29.764 20.826 ;
 END
 END vss.gds1821
 PIN vss.gds1822
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.474 21.6235 30.53 21.8235 ;
 END
 END vss.gds1822
 PIN vss.gds1823
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.646 25.031 33.702 25.231 ;
 END
 END vss.gds1823
 PIN vss.gds1824
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 23.2245 33.198 23.4245 ;
 END
 END vss.gds1824
 PIN vss.gds1825
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 24.37 34.366 24.57 ;
 END
 END vss.gds1825
 PIN vss.gds1826
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.65 23.595 34.706 23.795 ;
 END
 END vss.gds1826
 PIN vss.gds1827
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.314 21.568 31.37 21.768 ;
 END
 END vss.gds1827
 PIN vss.gds1828
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 21.779 31.922 21.979 ;
 END
 END vss.gds1828
 PIN vss.gds1829
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 23.1285 32.214 23.3285 ;
 END
 END vss.gds1829
 PIN vss.gds1830
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.222 24.6335 33.278 24.8335 ;
 END
 END vss.gds1830
 PIN vss.gds1831
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 23.2295 34.046 23.4295 ;
 END
 END vss.gds1831
 PIN vss.gds1832
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 23.041 30.71 23.241 ;
 END
 END vss.gds1832
 PIN vss.gds1833
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 23.427 32.894 23.627 ;
 END
 END vss.gds1833
 PIN vss.gds1834
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 23.128 33.542 23.328 ;
 END
 END vss.gds1834
 PIN vss.gds1835
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 23.111 31.55 23.311 ;
 END
 END vss.gds1835
 PIN vss.gds1836
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 21.426 33.866 21.626 ;
 END
 END vss.gds1836
 PIN vss.gds1837
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 23.2755 34.886 23.4755 ;
 END
 END vss.gds1837
 PIN vss.gds1838
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 21.568 32.47 21.768 ;
 END
 END vss.gds1838
 PIN vss.gds1839
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 20.957 34.366 21.157 ;
 END
 END vss.gds1839
 PIN vss.gds1840
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 31.304 24.759 31.36 24.941 ;
 RECT 32.144 24.819 32.2 25.019 ;
 RECT 31.808 24.778 31.864 24.978 ;
 RECT 31.556 24.759 31.612 24.941 ;
 RECT 32.48 24.778 32.536 24.978 ;
 RECT 33.068 24.778 33.124 24.978 ;
 RECT 32.9 24.778 32.956 24.978 ;
 RECT 33.572 24.759 33.628 24.941 ;
 RECT 33.32 24.759 33.376 24.941 ;
 RECT 34.16 24.778 34.216 24.978 ;
 RECT 34.328 24.778 34.384 24.978 ;
 RECT 30.296 22.071 30.352 22.253 ;
 RECT 32.984 22.09 33.04 22.29 ;
 RECT 32.816 22.09 32.872 22.29 ;
 RECT 32.648 22.09 32.704 22.29 ;
 RECT 32.48 22.09 32.536 22.29 ;
 RECT 33.656 22.09 33.712 22.29 ;
 RECT 33.236 22.072 33.292 22.249 ;
 RECT 30.296 21.847 30.352 22.029 ;
 RECT 30.968 21.95 31.024 22.15 ;
 RECT 32.984 21.81 33.04 22.01 ;
 RECT 32.816 21.81 32.872 22.01 ;
 RECT 32.648 21.81 32.704 22.01 ;
 RECT 32.48 21.81 32.536 22.01 ;
 RECT 33.236 21.851 33.292 22.029 ;
 RECT 33.404 21.847 33.46 22.047 ;
 RECT 33.74 21.81 33.796 22.01 ;
 RECT 34.916 21.81 34.972 22.01 ;
 RECT 30.548 23.154 30.604 23.354 ;
 RECT 30.968 23.154 31.024 23.354 ;
 RECT 31.388 23.154 31.444 23.354 ;
 RECT 31.892 23.154 31.948 23.354 ;
 RECT 31.724 23.191 31.78 23.373 ;
 RECT 32.228 23.0835 32.284 23.2835 ;
 RECT 33.152 23.195 33.208 23.367 ;
 RECT 32.9 23.195 32.956 23.367 ;
 RECT 32.564 23.154 32.62 23.354 ;
 RECT 33.572 23.154 33.628 23.354 ;
 RECT 34.58 23.154 34.636 23.354 ;
 RECT 34.076 23.154 34.132 23.354 ;
 RECT 31.724 23.415 31.78 23.597 ;
 RECT 31.892 23.434 31.948 23.634 ;
 RECT 33.152 23.415 33.208 23.593 ;
 RECT 32.564 23.434 32.62 23.634 ;
 RECT 32.9 23.415 32.956 23.593 ;
 RECT 33.656 23.434 33.712 23.634 ;
 RECT 34.16 23.434 34.216 23.634 ;
 RECT 34.58 23.434 34.636 23.634 ;
 RECT 30.632 20.748 30.688 20.948 ;
 RECT 30.968 20.748 31.024 20.948 ;
 RECT 31.304 20.748 31.36 20.948 ;
 RECT 31.64 20.748 31.696 20.948 ;
 RECT 31.976 20.748 32.032 20.948 ;
 RECT 32.984 20.748 33.04 20.948 ;
 RECT 33.32 20.748 33.376 20.948 ;
 RECT 33.656 20.748 33.712 20.948 ;
 RECT 33.992 20.748 34.048 20.948 ;
 RECT 33.572 20.516 33.628 20.669 ;
 RECT 31.052 20.496 31.108 20.669 ;
 RECT 31.22 20.469 31.276 20.669 ;
 RECT 32.816 20.513 32.872 20.678 ;
 RECT 32.648 20.513 32.704 20.678 ;
 RECT 31.892 20.513 31.948 20.678 ;
 RECT 31.724 20.513 31.78 20.678 ;
 RECT 34.16 21.95 34.216 22.15 ;
 RECT 33.992 21.95 34.048 22.15 ;
 RECT 34.328 21.95 34.384 22.15 ;
 RECT 30.296 20.709 30.352 20.909 ;
 RECT 34.832 24.8485 34.888 25.0485 ;
 RECT 30.548 23.5045 30.604 23.7045 ;
 RECT 30.968 23.5045 31.024 23.7045 ;
 RECT 31.388 23.5045 31.444 23.7045 ;
 RECT 32.228 23.5045 32.284 23.7045 ;
 RECT 34.58 22.0615 34.636 22.2615 ;
 RECT 34.832 22.131 34.888 22.331 ;
 RECT 30.296 24.638 30.352 24.838 ;
 RECT 31.304 24.535 31.36 24.717 ;
 RECT 30.968 24.638 31.024 24.838 ;
 RECT 32.144 24.498 32.2 24.698 ;
 RECT 31.808 24.498 31.864 24.698 ;
 RECT 31.64 24.535 31.696 24.717 ;
 RECT 33.152 24.535 33.208 24.717 ;
 RECT 32.48 24.498 32.536 24.698 ;
 RECT 32.816 24.535 32.872 24.717 ;
 RECT 33.656 24.498 33.712 24.698 ;
 RECT 34.244 24.535 34.3 24.717 ;
 RECT 34.328 20.709 34.384 20.909 ;
 RECT 30.38 20.543 30.436 20.743 ;
 RECT 32.228 20.554 32.284 20.754 ;
 RECT 34.916 20.543 34.972 20.743 ;
 RECT 34.748 20.543 34.804 20.743 ;
 RECT 34.58 20.543 34.636 20.743 ;
 RECT 34.412 20.543 34.468 20.743 ;
 RECT 34.244 20.543 34.3 20.743 ;
 RECT 35.084 20.543 35.14 20.743 ;
 RECT 34.076 20.554 34.132 20.754 ;
 END
 END vss.gds1840
 PIN vss.gds1841
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.634 22.185 39.674 22.385 ;
 END
 END vss.gds1841
 PIN vss.gds1842
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.962 22.185 39.002 22.385 ;
 END
 END vss.gds1842
 PIN vss.gds1843
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.29 22.185 38.33 22.385 ;
 END
 END vss.gds1843
 PIN vss.gds1844
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.618 22.185 37.658 22.385 ;
 END
 END vss.gds1844
 PIN vss.gds1845
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.946 22.185 36.986 22.385 ;
 END
 END vss.gds1845
 PIN vss.gds1846
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.274 22.185 36.314 22.385 ;
 END
 END vss.gds1846
 PIN vss.gds1847
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.102 22.49 40.148 22.69 ;
 END
 END vss.gds1847
 PIN vss.gds1848
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.43 22.49 39.476 22.69 ;
 END
 END vss.gds1848
 PIN vss.gds1849
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.826 22.6675 39.866 22.8675 ;
 END
 END vss.gds1849
 PIN vss.gds1850
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.758 22.49 38.804 22.69 ;
 END
 END vss.gds1850
 PIN vss.gds1851
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.154 22.6675 39.194 22.8675 ;
 END
 END vss.gds1851
 PIN vss.gds1852
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.086 22.49 38.132 22.69 ;
 END
 END vss.gds1852
 PIN vss.gds1853
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.482 22.6675 38.522 22.8675 ;
 END
 END vss.gds1853
 PIN vss.gds1854
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.414 22.49 37.46 22.69 ;
 END
 END vss.gds1854
 PIN vss.gds1855
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.81 22.6675 37.85 22.8675 ;
 END
 END vss.gds1855
 PIN vss.gds1856
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.742 22.49 36.788 22.69 ;
 END
 END vss.gds1856
 PIN vss.gds1857
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.138 22.6675 37.178 22.8675 ;
 END
 END vss.gds1857
 PIN vss.gds1858
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.07 22.49 36.116 22.69 ;
 END
 END vss.gds1858
 PIN vss.gds1859
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.466 22.6675 36.506 22.8675 ;
 END
 END vss.gds1859
 PIN vss.gds1860
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.398 22.49 35.444 22.69 ;
 END
 END vss.gds1860
 PIN vss.gds1861
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.794 22.6675 35.834 22.8675 ;
 END
 END vss.gds1861
 PIN vss.gds1862
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 23.1945 36.654 23.3945 ;
 END
 END vss.gds1862
 PIN vss.gds1863
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 23.1945 37.326 23.3945 ;
 END
 END vss.gds1863
 PIN vss.gds1864
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 23.1945 37.998 23.3945 ;
 END
 END vss.gds1864
 PIN vss.gds1865
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.602 22.185 35.642 22.385 ;
 END
 END vss.gds1865
 PIN vss.gds1866
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 23.1945 38.67 23.3945 ;
 END
 END vss.gds1866
 PIN vss.gds1867
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 23.1945 35.982 23.3945 ;
 END
 END vss.gds1867
 PIN vss.gds1868
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 23.1945 40.014 23.3945 ;
 END
 END vss.gds1868
 PIN vss.gds1869
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 23.1945 35.31 23.3945 ;
 END
 END vss.gds1869
 PIN vss.gds1870
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 23.1945 39.342 23.3945 ;
 END
 END vss.gds1870
 PIN vss.gds1871
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 35.252 24.302 35.308 24.502 ;
 RECT 40.124 22.7325 40.18 22.9325 ;
 RECT 39.62 22.7325 39.676 22.9325 ;
 RECT 39.452 22.7325 39.508 22.9325 ;
 RECT 39.956 22.7325 40.012 22.9325 ;
 RECT 39.788 22.7325 39.844 22.9325 ;
 RECT 38.948 22.7325 39.004 22.9325 ;
 RECT 38.78 22.7325 38.836 22.9325 ;
 RECT 39.284 22.7325 39.34 22.9325 ;
 RECT 39.116 22.7325 39.172 22.9325 ;
 RECT 38.276 22.7325 38.332 22.9325 ;
 RECT 38.108 22.7325 38.164 22.9325 ;
 RECT 38.612 22.7325 38.668 22.9325 ;
 RECT 38.444 22.7325 38.5 22.9325 ;
 RECT 37.604 22.7325 37.66 22.9325 ;
 RECT 37.436 22.7325 37.492 22.9325 ;
 RECT 37.94 22.7325 37.996 22.9325 ;
 RECT 37.772 22.7325 37.828 22.9325 ;
 RECT 36.932 22.7325 36.988 22.9325 ;
 RECT 36.764 22.7325 36.82 22.9325 ;
 RECT 37.268 22.7325 37.324 22.9325 ;
 RECT 37.1 22.7325 37.156 22.9325 ;
 RECT 36.26 22.7325 36.316 22.9325 ;
 RECT 36.092 22.7325 36.148 22.9325 ;
 RECT 36.596 22.7325 36.652 22.9325 ;
 RECT 36.428 22.7325 36.484 22.9325 ;
 RECT 35.588 22.7325 35.644 22.9325 ;
 RECT 35.252 22.7325 35.308 22.9325 ;
 RECT 35.42 22.7325 35.476 22.9325 ;
 RECT 35.924 22.7325 35.98 22.9325 ;
 RECT 35.756 22.7325 35.812 22.9325 ;
 RECT 39.956 24.5075 40.012 24.7075 ;
 RECT 39.284 24.5075 39.34 24.7075 ;
 RECT 38.612 24.5075 38.668 24.7075 ;
 RECT 37.94 24.5075 37.996 24.7075 ;
 RECT 37.268 24.5075 37.324 24.7075 ;
 RECT 36.596 24.5075 36.652 24.7075 ;
 RECT 35.924 24.5075 35.98 24.7075 ;
 RECT 40.124 21.19 40.18 21.39 ;
 RECT 39.62 21.19 39.676 21.39 ;
 RECT 39.452 21.19 39.508 21.39 ;
 RECT 39.788 21.19 39.844 21.39 ;
 RECT 39.956 21.181 40.012 21.381 ;
 RECT 38.948 21.19 39.004 21.39 ;
 RECT 38.78 21.19 38.836 21.39 ;
 RECT 39.116 21.19 39.172 21.39 ;
 RECT 39.284 21.181 39.34 21.381 ;
 RECT 38.276 21.19 38.332 21.39 ;
 RECT 38.108 21.19 38.164 21.39 ;
 RECT 38.444 21.19 38.5 21.39 ;
 RECT 38.612 21.181 38.668 21.381 ;
 RECT 37.604 21.19 37.66 21.39 ;
 RECT 37.436 21.19 37.492 21.39 ;
 RECT 37.772 21.19 37.828 21.39 ;
 RECT 37.94 21.181 37.996 21.381 ;
 RECT 36.932 21.19 36.988 21.39 ;
 RECT 36.764 21.19 36.82 21.39 ;
 RECT 37.1 21.19 37.156 21.39 ;
 RECT 37.268 21.181 37.324 21.381 ;
 RECT 36.26 21.19 36.316 21.39 ;
 RECT 36.092 21.19 36.148 21.39 ;
 RECT 36.428 21.19 36.484 21.39 ;
 RECT 36.596 21.181 36.652 21.381 ;
 RECT 35.252 21.181 35.308 21.381 ;
 RECT 35.588 21.19 35.644 21.39 ;
 RECT 35.42 21.19 35.476 21.39 ;
 RECT 35.756 21.19 35.812 21.39 ;
 RECT 35.924 21.181 35.98 21.381 ;
 END
 END vss.gds1871
 PIN vss.gds1872
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.758 22.185 44.798 22.385 ;
 END
 END vss.gds1872
 PIN vss.gds1873
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.086 22.185 44.126 22.385 ;
 END
 END vss.gds1873
 PIN vss.gds1874
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.414 22.185 43.454 22.385 ;
 END
 END vss.gds1874
 PIN vss.gds1875
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.742 22.185 42.782 22.385 ;
 END
 END vss.gds1875
 PIN vss.gds1876
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.07 22.185 42.11 22.385 ;
 END
 END vss.gds1876
 PIN vss.gds1877
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.398 22.185 41.438 22.385 ;
 END
 END vss.gds1877
 PIN vss.gds1878
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.306 22.185 40.346 22.385 ;
 END
 END vss.gds1878
 PIN vss.gds1879
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.226 22.49 45.272 22.69 ;
 END
 END vss.gds1879
 PIN vss.gds1880
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.554 22.49 44.6 22.69 ;
 END
 END vss.gds1880
 PIN vss.gds1881
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.95 22.6675 44.99 22.8675 ;
 END
 END vss.gds1881
 PIN vss.gds1882
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.882 22.49 43.928 22.69 ;
 END
 END vss.gds1882
 PIN vss.gds1883
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.278 22.6675 44.318 22.8675 ;
 END
 END vss.gds1883
 PIN vss.gds1884
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.21 22.49 43.256 22.69 ;
 END
 END vss.gds1884
 PIN vss.gds1885
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.606 22.6675 43.646 22.8675 ;
 END
 END vss.gds1885
 PIN vss.gds1886
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.538 22.49 42.584 22.69 ;
 END
 END vss.gds1886
 PIN vss.gds1887
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.934 22.6675 42.974 22.8675 ;
 END
 END vss.gds1887
 PIN vss.gds1888
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.866 22.49 41.912 22.69 ;
 END
 END vss.gds1888
 PIN vss.gds1889
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.262 22.6675 42.302 22.8675 ;
 END
 END vss.gds1889
 PIN vss.gds1890
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.194 22.49 41.24 22.69 ;
 END
 END vss.gds1890
 PIN vss.gds1891
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.59 22.6675 41.63 22.8675 ;
 END
 END vss.gds1891
 PIN vss.gds1892
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.498 22.6675 40.538 22.8675 ;
 END
 END vss.gds1892
 PIN vss.gds1893
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.774 23.932 40.814 24.132 ;
 END
 END vss.gds1893
 PIN vss.gds1894
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.918 23.932 40.958 24.132 ;
 END
 END vss.gds1894
 PIN vss.gds1895
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 23.1945 45.138 23.3945 ;
 END
 END vss.gds1895
 PIN vss.gds1896
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 23.1945 44.466 23.3945 ;
 END
 END vss.gds1896
 PIN vss.gds1897
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 23.1945 43.794 23.3945 ;
 END
 END vss.gds1897
 PIN vss.gds1898
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 23.1945 43.122 23.3945 ;
 END
 END vss.gds1898
 PIN vss.gds1899
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 23.1945 42.45 23.3945 ;
 END
 END vss.gds1899
 PIN vss.gds1900
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 23.1945 41.778 23.3945 ;
 END
 END vss.gds1900
 PIN vss.gds1901
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 23.2565 40.686 23.4565 ;
 END
 END vss.gds1901
 PIN vss.gds1902
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.046 23.2565 41.106 23.4565 ;
 END
 END vss.gds1902
 PIN vss.gds1903
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 44.744 21.19 44.8 21.39 ;
 RECT 44.576 21.19 44.632 21.39 ;
 RECT 44.912 21.19 44.968 21.39 ;
 RECT 45.08 21.181 45.136 21.381 ;
 RECT 44.072 21.19 44.128 21.39 ;
 RECT 43.904 21.19 43.96 21.39 ;
 RECT 44.24 21.19 44.296 21.39 ;
 RECT 44.408 21.181 44.464 21.381 ;
 RECT 43.4 21.19 43.456 21.39 ;
 RECT 43.232 21.19 43.288 21.39 ;
 RECT 43.568 21.19 43.624 21.39 ;
 RECT 43.736 21.181 43.792 21.381 ;
 RECT 42.728 21.19 42.784 21.39 ;
 RECT 42.56 21.19 42.616 21.39 ;
 RECT 42.896 21.19 42.952 21.39 ;
 RECT 43.064 21.181 43.12 21.381 ;
 RECT 42.056 21.19 42.112 21.39 ;
 RECT 41.888 21.19 41.944 21.39 ;
 RECT 42.224 21.19 42.28 21.39 ;
 RECT 42.392 21.181 42.448 21.381 ;
 RECT 41.72 21.181 41.776 21.381 ;
 RECT 40.628 21.181 40.684 21.381 ;
 RECT 41.048 21.0105 41.104 21.2105 ;
 RECT 41.384 21.19 41.44 21.39 ;
 RECT 41.216 21.19 41.272 21.39 ;
 RECT 41.552 21.19 41.608 21.39 ;
 RECT 41.048 24.302 41.104 24.502 ;
 RECT 44.744 22.7325 44.8 22.9325 ;
 RECT 44.576 22.7325 44.632 22.9325 ;
 RECT 45.08 22.7325 45.136 22.9325 ;
 RECT 44.912 22.7325 44.968 22.9325 ;
 RECT 44.072 22.7325 44.128 22.9325 ;
 RECT 43.904 22.7325 43.96 22.9325 ;
 RECT 44.408 22.7325 44.464 22.9325 ;
 RECT 44.24 22.7325 44.296 22.9325 ;
 RECT 43.4 22.7325 43.456 22.9325 ;
 RECT 43.232 22.7325 43.288 22.9325 ;
 RECT 43.736 22.7325 43.792 22.9325 ;
 RECT 43.568 22.7325 43.624 22.9325 ;
 RECT 42.728 22.7325 42.784 22.9325 ;
 RECT 42.56 22.7325 42.616 22.9325 ;
 RECT 43.064 22.7325 43.12 22.9325 ;
 RECT 42.896 22.7325 42.952 22.9325 ;
 RECT 42.056 22.7325 42.112 22.9325 ;
 RECT 41.888 22.7325 41.944 22.9325 ;
 RECT 42.392 22.7325 42.448 22.9325 ;
 RECT 42.224 22.7325 42.28 22.9325 ;
 RECT 41.384 22.7325 41.44 22.9325 ;
 RECT 41.048 22.7325 41.104 22.9325 ;
 RECT 41.216 22.7325 41.272 22.9325 ;
 RECT 41.72 22.7325 41.776 22.9325 ;
 RECT 41.552 22.7325 41.608 22.9325 ;
 RECT 40.628 22.7325 40.684 22.9325 ;
 RECT 40.46 22.7325 40.516 22.9325 ;
 RECT 40.292 22.7325 40.348 22.9325 ;
 RECT 45.08 24.5075 45.136 24.7075 ;
 RECT 44.408 24.5075 44.464 24.7075 ;
 RECT 43.736 24.5075 43.792 24.7075 ;
 RECT 43.064 24.5075 43.12 24.7075 ;
 RECT 42.392 24.5075 42.448 24.7075 ;
 RECT 41.72 24.5075 41.776 24.7075 ;
 RECT 40.628 24.5075 40.684 24.7075 ;
 RECT 40.46 21.19 40.516 21.39 ;
 RECT 40.292 21.19 40.348 21.39 ;
 RECT 40.796 22.7795 40.852 22.9795 ;
 END
 END vss.gds1903
 PIN vss.gds1904
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.102 22.185 46.142 22.385 ;
 END
 END vss.gds1904
 PIN vss.gds1905
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.43 22.185 45.47 22.385 ;
 END
 END vss.gds1905
 PIN vss.gds1906
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.898 22.49 45.944 22.69 ;
 END
 END vss.gds1906
 PIN vss.gds1907
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.294 22.6675 46.334 22.8675 ;
 END
 END vss.gds1907
 PIN vss.gds1908
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.622 22.6675 45.662 22.8675 ;
 END
 END vss.gds1908
 PIN vss.gds1909
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.366 21.568 48.422 21.768 ;
 END
 END vss.gds1909
 PIN vss.gds1910
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 21.615 47.162 21.815 ;
 END
 END vss.gds1910
 PIN vss.gds1911
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 23.2245 50.25 23.4245 ;
 END
 END vss.gds1911
 PIN vss.gds1912
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 21.779 48.974 21.979 ;
 END
 END vss.gds1912
 PIN vss.gds1913
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.526 21.6235 47.582 21.8235 ;
 END
 END vss.gds1913
 PIN vss.gds1914
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 23.0545 46.482 23.2545 ;
 END
 END vss.gds1914
 PIN vss.gds1915
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 23.1945 45.81 23.3945 ;
 END
 END vss.gds1915
 PIN vss.gds1916
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 23.041 46.922 23.241 ;
 END
 END vss.gds1916
 PIN vss.gds1917
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 23.3375 46.694 23.5375 ;
 END
 END vss.gds1917
 PIN vss.gds1918
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 23.041 47.762 23.241 ;
 END
 END vss.gds1918
 PIN vss.gds1919
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 23.1285 49.266 23.3285 ;
 END
 END vss.gds1919
 PIN vss.gds1920
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 23.111 48.602 23.311 ;
 END
 END vss.gds1920
 PIN vss.gds1921
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 23.427 49.946 23.627 ;
 END
 END vss.gds1921
 PIN vss.gds1922
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 21.568 49.522 21.768 ;
 END
 END vss.gds1922
 PIN vss.gds1923
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 46.844 24.778 46.9 24.978 ;
 RECT 48.356 24.759 48.412 24.941 ;
 RECT 49.196 24.819 49.252 25.019 ;
 RECT 48.86 24.778 48.916 24.978 ;
 RECT 48.608 24.759 48.664 24.941 ;
 RECT 49.532 24.778 49.588 24.978 ;
 RECT 50.12 24.778 50.176 24.978 ;
 RECT 49.952 24.778 50.008 24.978 ;
 RECT 46.76 22.09 46.816 22.29 ;
 RECT 47.348 22.071 47.404 22.253 ;
 RECT 50.036 22.09 50.092 22.29 ;
 RECT 49.868 22.09 49.924 22.29 ;
 RECT 49.7 22.09 49.756 22.29 ;
 RECT 49.532 22.09 49.588 22.29 ;
 RECT 46.76 21.81 46.816 22.01 ;
 RECT 47.348 21.847 47.404 22.029 ;
 RECT 48.02 21.95 48.076 22.15 ;
 RECT 50.036 21.81 50.092 22.01 ;
 RECT 49.868 21.81 49.924 22.01 ;
 RECT 49.7 21.81 49.756 22.01 ;
 RECT 49.532 21.81 49.588 22.01 ;
 RECT 47.6 23.154 47.656 23.354 ;
 RECT 47.18 23.154 47.236 23.354 ;
 RECT 48.02 23.154 48.076 23.354 ;
 RECT 48.44 23.154 48.496 23.354 ;
 RECT 48.944 23.154 49 23.354 ;
 RECT 48.776 23.191 48.832 23.373 ;
 RECT 49.28 23.0835 49.336 23.2835 ;
 RECT 50.204 23.195 50.26 23.367 ;
 RECT 49.952 23.195 50.008 23.367 ;
 RECT 49.616 23.154 49.672 23.354 ;
 RECT 48.776 23.415 48.832 23.597 ;
 RECT 48.944 23.434 49 23.634 ;
 RECT 50.204 23.415 50.26 23.593 ;
 RECT 49.616 23.434 49.672 23.634 ;
 RECT 49.952 23.415 50.008 23.593 ;
 RECT 47.684 20.748 47.74 20.948 ;
 RECT 47.012 20.748 47.068 20.948 ;
 RECT 48.02 20.748 48.076 20.948 ;
 RECT 48.356 20.748 48.412 20.948 ;
 RECT 48.692 20.748 48.748 20.948 ;
 RECT 49.028 20.748 49.084 20.948 ;
 RECT 50.036 20.748 50.092 20.948 ;
 RECT 47.348 20.709 47.404 20.909 ;
 RECT 46.088 21.19 46.144 21.39 ;
 RECT 46.424 21.181 46.48 21.381 ;
 RECT 45.416 21.19 45.472 21.39 ;
 RECT 45.248 21.19 45.304 21.39 ;
 RECT 45.584 21.19 45.64 21.39 ;
 RECT 45.752 21.181 45.808 21.381 ;
 RECT 48.104 20.496 48.16 20.669 ;
 RECT 48.272 20.469 48.328 20.669 ;
 RECT 49.868 20.513 49.924 20.678 ;
 RECT 49.7 20.513 49.756 20.678 ;
 RECT 48.944 20.513 49 20.678 ;
 RECT 48.776 20.513 48.832 20.678 ;
 RECT 47.18 23.5045 47.236 23.7045 ;
 RECT 47.6 23.5045 47.656 23.7045 ;
 RECT 48.02 23.5045 48.076 23.7045 ;
 RECT 48.44 23.5045 48.496 23.7045 ;
 RECT 49.28 23.5045 49.336 23.7045 ;
 RECT 47.348 24.638 47.404 24.838 ;
 RECT 48.356 24.535 48.412 24.717 ;
 RECT 48.02 24.638 48.076 24.838 ;
 RECT 49.196 24.498 49.252 24.698 ;
 RECT 48.86 24.498 48.916 24.698 ;
 RECT 48.692 24.535 48.748 24.717 ;
 RECT 50.204 24.535 50.26 24.717 ;
 RECT 49.532 24.498 49.588 24.698 ;
 RECT 49.868 24.535 49.924 24.717 ;
 RECT 46.088 22.7325 46.144 22.9325 ;
 RECT 45.92 22.7325 45.976 22.9325 ;
 RECT 46.424 22.7325 46.48 22.9325 ;
 RECT 46.256 22.7325 46.312 22.9325 ;
 RECT 45.416 22.7325 45.472 22.9325 ;
 RECT 45.248 22.7325 45.304 22.9325 ;
 RECT 45.752 22.7325 45.808 22.9325 ;
 RECT 45.584 22.7325 45.64 22.9325 ;
 RECT 46.424 24.5075 46.48 24.7075 ;
 RECT 45.752 24.5075 45.808 24.7075 ;
 RECT 47.432 20.543 47.488 20.743 ;
 RECT 47.264 20.543 47.32 20.743 ;
 RECT 46.928 20.543 46.984 20.743 ;
 RECT 47.096 20.543 47.152 20.743 ;
 RECT 49.28 20.554 49.336 20.754 ;
 RECT 46.592 20.543 46.648 20.743 ;
 RECT 45.92 21.19 45.976 21.39 ;
 RECT 46.256 21.19 46.312 21.39 ;
 RECT 46.76 20.626 46.816 20.826 ;
 END
 END vss.gds1923
 PIN vss.gds1924
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.138 22.49 55.184 22.69 ;
 END
 END vss.gds1924
 PIN vss.gds1925
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.466 22.49 54.512 22.69 ;
 END
 END vss.gds1925
 PIN vss.gds1926
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.794 22.49 53.84 22.69 ;
 END
 END vss.gds1926
 PIN vss.gds1927
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.122 22.49 53.168 22.69 ;
 END
 END vss.gds1927
 PIN vss.gds1928
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.45 22.49 52.496 22.69 ;
 END
 END vss.gds1928
 PIN vss.gds1929
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.698 25.031 50.754 25.231 ;
 END
 END vss.gds1929
 PIN vss.gds1930
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.702 23.595 51.758 23.795 ;
 END
 END vss.gds1930
 PIN vss.gds1931
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.846 22.6675 52.886 22.8675 ;
 END
 END vss.gds1931
 PIN vss.gds1932
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.518 22.6675 53.558 22.8675 ;
 END
 END vss.gds1932
 PIN vss.gds1933
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.67 22.185 54.71 22.385 ;
 END
 END vss.gds1933
 PIN vss.gds1934
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 23.1945 55.05 23.3945 ;
 END
 END vss.gds1934
 PIN vss.gds1935
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 23.1945 54.378 23.3945 ;
 END
 END vss.gds1935
 PIN vss.gds1936
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.862 22.6675 54.902 22.8675 ;
 END
 END vss.gds1936
 PIN vss.gds1937
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.998 22.185 54.038 22.385 ;
 END
 END vss.gds1937
 PIN vss.gds1938
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.19 22.6675 54.23 22.8675 ;
 END
 END vss.gds1938
 PIN vss.gds1939
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.326 22.185 53.366 22.385 ;
 END
 END vss.gds1939
 PIN vss.gds1940
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.654 22.185 52.694 22.385 ;
 END
 END vss.gds1940
 PIN vss.gds1941
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 24.37 51.418 24.57 ;
 END
 END vss.gds1941
 PIN vss.gds1942
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 21.426 50.918 21.626 ;
 END
 END vss.gds1942
 PIN vss.gds1943
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 23.1945 53.706 23.3945 ;
 END
 END vss.gds1943
 PIN vss.gds1944
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.274 24.6335 50.33 24.8335 ;
 END
 END vss.gds1944
 PIN vss.gds1945
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 23.2295 51.098 23.4295 ;
 END
 END vss.gds1945
 PIN vss.gds1946
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 23.1945 53.034 23.3945 ;
 END
 END vss.gds1946
 PIN vss.gds1947
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 23.2755 51.938 23.4755 ;
 END
 END vss.gds1947
 PIN vss.gds1948
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 20.957 51.418 21.157 ;
 END
 END vss.gds1948
 PIN vss.gds1949
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 23.128 50.594 23.328 ;
 END
 END vss.gds1949
 PIN vss.gds1950
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 23.1945 52.362 23.3945 ;
 END
 END vss.gds1950
 PIN vss.gds1951
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 50.624 24.759 50.68 24.941 ;
 RECT 50.372 24.759 50.428 24.941 ;
 RECT 51.212 24.778 51.268 24.978 ;
 RECT 51.38 24.778 51.436 24.978 ;
 RECT 50.708 22.09 50.764 22.29 ;
 RECT 50.288 22.072 50.344 22.249 ;
 RECT 50.288 21.851 50.344 22.029 ;
 RECT 50.456 21.847 50.512 22.047 ;
 RECT 50.792 21.81 50.848 22.01 ;
 RECT 51.968 21.81 52.024 22.01 ;
 RECT 50.624 23.154 50.68 23.354 ;
 RECT 51.632 23.154 51.688 23.354 ;
 RECT 51.128 23.154 51.184 23.354 ;
 RECT 50.708 23.434 50.764 23.634 ;
 RECT 51.212 23.434 51.268 23.634 ;
 RECT 51.632 23.434 51.688 23.634 ;
 RECT 50.372 20.748 50.428 20.948 ;
 RECT 50.708 20.748 50.764 20.948 ;
 RECT 51.044 20.748 51.1 20.948 ;
 RECT 50.624 20.516 50.68 20.669 ;
 RECT 55.16 22.7325 55.216 22.9325 ;
 RECT 54.656 22.7325 54.712 22.9325 ;
 RECT 54.488 22.7325 54.544 22.9325 ;
 RECT 54.992 22.7325 55.048 22.9325 ;
 RECT 54.824 22.7325 54.88 22.9325 ;
 RECT 53.984 22.7325 54.04 22.9325 ;
 RECT 53.816 22.7325 53.872 22.9325 ;
 RECT 54.32 22.7325 54.376 22.9325 ;
 RECT 54.152 22.7325 54.208 22.9325 ;
 RECT 53.312 22.7325 53.368 22.9325 ;
 RECT 53.144 22.7325 53.2 22.9325 ;
 RECT 53.648 22.7325 53.704 22.9325 ;
 RECT 53.48 22.7325 53.536 22.9325 ;
 RECT 52.64 22.7325 52.696 22.9325 ;
 RECT 52.304 22.7325 52.36 22.9325 ;
 RECT 52.472 22.7325 52.528 22.9325 ;
 RECT 52.976 22.7325 53.032 22.9325 ;
 RECT 52.808 22.7325 52.864 22.9325 ;
 RECT 51.212 21.95 51.268 22.15 ;
 RECT 51.044 21.95 51.1 22.15 ;
 RECT 51.38 21.95 51.436 22.15 ;
 RECT 51.884 24.8485 51.94 25.0485 ;
 RECT 51.632 22.0615 51.688 22.2615 ;
 RECT 51.884 22.131 51.94 22.331 ;
 RECT 54.992 24.5075 55.048 24.7075 ;
 RECT 54.32 24.5075 54.376 24.7075 ;
 RECT 53.648 24.5075 53.704 24.7075 ;
 RECT 52.304 24.302 52.36 24.502 ;
 RECT 52.976 24.5075 53.032 24.7075 ;
 RECT 50.708 24.498 50.764 24.698 ;
 RECT 51.296 24.535 51.352 24.717 ;
 RECT 55.16 21.19 55.216 21.39 ;
 RECT 54.656 21.19 54.712 21.39 ;
 RECT 54.488 21.19 54.544 21.39 ;
 RECT 54.824 21.19 54.88 21.39 ;
 RECT 54.992 21.181 55.048 21.381 ;
 RECT 53.984 21.19 54.04 21.39 ;
 RECT 53.816 21.19 53.872 21.39 ;
 RECT 54.152 21.19 54.208 21.39 ;
 RECT 54.32 21.181 54.376 21.381 ;
 RECT 53.312 21.19 53.368 21.39 ;
 RECT 53.144 21.19 53.2 21.39 ;
 RECT 53.48 21.19 53.536 21.39 ;
 RECT 53.648 21.181 53.704 21.381 ;
 RECT 52.304 21.181 52.36 21.381 ;
 RECT 51.38 20.709 51.436 20.909 ;
 RECT 52.64 21.19 52.696 21.39 ;
 RECT 52.472 21.19 52.528 21.39 ;
 RECT 52.808 21.19 52.864 21.39 ;
 RECT 52.976 21.181 53.032 21.381 ;
 RECT 51.968 20.543 52.024 20.743 ;
 RECT 51.8 20.543 51.856 20.743 ;
 RECT 51.632 20.543 51.688 20.743 ;
 RECT 51.464 20.543 51.52 20.743 ;
 RECT 51.296 20.543 51.352 20.743 ;
 RECT 52.136 20.543 52.192 20.743 ;
 RECT 51.128 20.554 51.184 20.754 ;
 END
 END vss.gds1951
 PIN vss.gds1952
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.59 22.49 59.636 22.69 ;
 END
 END vss.gds1952
 PIN vss.gds1953
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.918 22.49 58.964 22.69 ;
 END
 END vss.gds1953
 PIN vss.gds1954
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.246 22.49 58.292 22.69 ;
 END
 END vss.gds1954
 PIN vss.gds1955
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.154 22.49 57.2 22.69 ;
 END
 END vss.gds1955
 PIN vss.gds1956
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.482 22.49 56.528 22.69 ;
 END
 END vss.gds1956
 PIN vss.gds1957
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.81 22.49 55.856 22.69 ;
 END
 END vss.gds1957
 PIN vss.gds1958
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.826 23.932 57.866 24.132 ;
 END
 END vss.gds1958
 PIN vss.gds1959
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.97 23.932 58.01 24.132 ;
 END
 END vss.gds1959
 PIN vss.gds1960
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.794 22.185 59.834 22.385 ;
 END
 END vss.gds1960
 PIN vss.gds1961
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.986 22.6675 60.026 22.8675 ;
 END
 END vss.gds1961
 PIN vss.gds1962
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.122 22.185 59.162 22.385 ;
 END
 END vss.gds1962
 PIN vss.gds1963
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.314 22.6675 59.354 22.8675 ;
 END
 END vss.gds1963
 PIN vss.gds1964
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.45 22.185 58.49 22.385 ;
 END
 END vss.gds1964
 PIN vss.gds1965
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.642 22.6675 58.682 22.8675 ;
 END
 END vss.gds1965
 PIN vss.gds1966
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.358 22.185 57.398 22.385 ;
 END
 END vss.gds1966
 PIN vss.gds1967
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.55 22.6675 57.59 22.8675 ;
 END
 END vss.gds1967
 PIN vss.gds1968
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.686 22.185 56.726 22.385 ;
 END
 END vss.gds1968
 PIN vss.gds1969
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.878 22.6675 56.918 22.8675 ;
 END
 END vss.gds1969
 PIN vss.gds1970
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.014 22.185 56.054 22.385 ;
 END
 END vss.gds1970
 PIN vss.gds1971
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.206 22.6675 56.246 22.8675 ;
 END
 END vss.gds1971
 PIN vss.gds1972
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.342 22.185 55.382 22.385 ;
 END
 END vss.gds1972
 PIN vss.gds1973
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.534 22.6675 55.574 22.8675 ;
 END
 END vss.gds1973
 PIN vss.gds1974
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.098 23.2565 58.158 23.4565 ;
 END
 END vss.gds1974
 PIN vss.gds1975
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 23.1945 60.174 23.3945 ;
 END
 END vss.gds1975
 PIN vss.gds1976
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 23.1945 59.502 23.3945 ;
 END
 END vss.gds1976
 PIN vss.gds1977
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 23.1945 58.83 23.3945 ;
 END
 END vss.gds1977
 PIN vss.gds1978
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 23.1945 55.722 23.3945 ;
 END
 END vss.gds1978
 PIN vss.gds1979
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 23.1945 56.394 23.3945 ;
 END
 END vss.gds1979
 PIN vss.gds1980
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 23.2565 57.738 23.4565 ;
 END
 END vss.gds1980
 PIN vss.gds1981
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 23.1945 57.066 23.3945 ;
 END
 END vss.gds1981
 PIN vss.gds1982
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 59.78 22.7325 59.836 22.9325 ;
 RECT 59.612 22.7325 59.668 22.9325 ;
 RECT 60.116 22.7325 60.172 22.9325 ;
 RECT 59.948 22.7325 60.004 22.9325 ;
 RECT 59.108 22.7325 59.164 22.9325 ;
 RECT 58.94 22.7325 58.996 22.9325 ;
 RECT 59.444 22.7325 59.5 22.9325 ;
 RECT 59.276 22.7325 59.332 22.9325 ;
 RECT 58.436 22.7325 58.492 22.9325 ;
 RECT 58.1 22.7325 58.156 22.9325 ;
 RECT 58.268 22.7325 58.324 22.9325 ;
 RECT 58.772 22.7325 58.828 22.9325 ;
 RECT 58.604 22.7325 58.66 22.9325 ;
 RECT 57.344 22.7325 57.4 22.9325 ;
 RECT 57.176 22.7325 57.232 22.9325 ;
 RECT 57.68 22.7325 57.736 22.9325 ;
 RECT 57.512 22.7325 57.568 22.9325 ;
 RECT 56.672 22.7325 56.728 22.9325 ;
 RECT 56.504 22.7325 56.56 22.9325 ;
 RECT 57.008 22.7325 57.064 22.9325 ;
 RECT 56.84 22.7325 56.896 22.9325 ;
 RECT 56 22.7325 56.056 22.9325 ;
 RECT 55.832 22.7325 55.888 22.9325 ;
 RECT 56.336 22.7325 56.392 22.9325 ;
 RECT 56.168 22.7325 56.224 22.9325 ;
 RECT 55.328 22.7325 55.384 22.9325 ;
 RECT 55.664 22.7325 55.72 22.9325 ;
 RECT 55.496 22.7325 55.552 22.9325 ;
 RECT 60.116 24.5075 60.172 24.7075 ;
 RECT 59.444 24.5075 59.5 24.7075 ;
 RECT 58.1 24.302 58.156 24.502 ;
 RECT 58.772 24.5075 58.828 24.7075 ;
 RECT 57.68 24.5075 57.736 24.7075 ;
 RECT 57.008 24.5075 57.064 24.7075 ;
 RECT 56.336 24.5075 56.392 24.7075 ;
 RECT 55.664 24.5075 55.72 24.7075 ;
 RECT 59.78 21.19 59.836 21.39 ;
 RECT 59.612 21.19 59.668 21.39 ;
 RECT 59.948 21.19 60.004 21.39 ;
 RECT 60.116 21.181 60.172 21.381 ;
 RECT 59.108 21.19 59.164 21.39 ;
 RECT 58.94 21.19 58.996 21.39 ;
 RECT 59.276 21.19 59.332 21.39 ;
 RECT 59.444 21.181 59.5 21.381 ;
 RECT 58.772 21.181 58.828 21.381 ;
 RECT 58.1 21.0105 58.156 21.2105 ;
 RECT 58.436 21.19 58.492 21.39 ;
 RECT 58.268 21.19 58.324 21.39 ;
 RECT 58.604 21.19 58.66 21.39 ;
 RECT 57.344 21.19 57.4 21.39 ;
 RECT 57.176 21.19 57.232 21.39 ;
 RECT 57.512 21.19 57.568 21.39 ;
 RECT 57.68 21.181 57.736 21.381 ;
 RECT 56.672 21.19 56.728 21.39 ;
 RECT 56.504 21.19 56.56 21.39 ;
 RECT 56.84 21.19 56.896 21.39 ;
 RECT 57.008 21.181 57.064 21.381 ;
 RECT 56 21.19 56.056 21.39 ;
 RECT 55.832 21.19 55.888 21.39 ;
 RECT 56.168 21.19 56.224 21.39 ;
 RECT 56.336 21.181 56.392 21.381 ;
 RECT 55.328 21.19 55.384 21.39 ;
 RECT 55.496 21.19 55.552 21.39 ;
 RECT 55.664 21.181 55.72 21.381 ;
 RECT 57.848 22.7795 57.904 22.9795 ;
 END
 END vss.gds1982
 PIN vss.gds1983
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.95 22.49 62.996 22.69 ;
 END
 END vss.gds1983
 PIN vss.gds1984
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.278 22.49 62.324 22.69 ;
 END
 END vss.gds1984
 PIN vss.gds1985
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.606 22.49 61.652 22.69 ;
 END
 END vss.gds1985
 PIN vss.gds1986
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.934 22.49 60.98 22.69 ;
 END
 END vss.gds1986
 PIN vss.gds1987
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.262 22.49 60.308 22.69 ;
 END
 END vss.gds1987
 PIN vss.gds1988
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 21.615 64.214 21.815 ;
 END
 END vss.gds1988
 PIN vss.gds1989
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.578 21.6235 64.634 21.8235 ;
 END
 END vss.gds1989
 PIN vss.gds1990
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.154 22.185 63.194 22.385 ;
 END
 END vss.gds1990
 PIN vss.gds1991
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.346 22.6675 63.386 22.8675 ;
 END
 END vss.gds1991
 PIN vss.gds1992
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.482 22.185 62.522 22.385 ;
 END
 END vss.gds1992
 PIN vss.gds1993
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.674 22.6675 62.714 22.8675 ;
 END
 END vss.gds1993
 PIN vss.gds1994
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.81 22.185 61.85 22.385 ;
 END
 END vss.gds1994
 PIN vss.gds1995
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.002 22.6675 62.042 22.8675 ;
 END
 END vss.gds1995
 PIN vss.gds1996
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.138 22.185 61.178 22.385 ;
 END
 END vss.gds1996
 PIN vss.gds1997
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.33 22.6675 61.37 22.8675 ;
 END
 END vss.gds1997
 PIN vss.gds1998
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.466 22.185 60.506 22.385 ;
 END
 END vss.gds1998
 PIN vss.gds1999
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.658 22.6675 60.698 22.8675 ;
 END
 END vss.gds1999
 PIN vss.gds2000
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 23.0545 63.534 23.2545 ;
 END
 END vss.gds2000
 PIN vss.gds2001
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 23.1945 62.862 23.3945 ;
 END
 END vss.gds2001
 PIN vss.gds2002
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 23.1945 62.19 23.3945 ;
 END
 END vss.gds2002
 PIN vss.gds2003
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 23.1945 61.518 23.3945 ;
 END
 END vss.gds2003
 PIN vss.gds2004
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 23.1945 60.846 23.3945 ;
 END
 END vss.gds2004
 PIN vss.gds2005
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 23.041 63.974 23.241 ;
 END
 END vss.gds2005
 PIN vss.gds2006
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 23.3375 63.746 23.5375 ;
 END
 END vss.gds2006
 PIN vss.gds2007
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 23.041 64.814 23.241 ;
 END
 END vss.gds2007
 PIN vss.gds2008
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 63.896 24.778 63.952 24.978 ;
 RECT 63.812 22.09 63.868 22.29 ;
 RECT 64.4 22.071 64.456 22.253 ;
 RECT 63.812 21.81 63.868 22.01 ;
 RECT 64.4 21.847 64.456 22.029 ;
 RECT 65.072 21.95 65.128 22.15 ;
 RECT 64.652 23.154 64.708 23.354 ;
 RECT 64.232 23.154 64.288 23.354 ;
 RECT 65.072 23.154 65.128 23.354 ;
 RECT 64.736 20.748 64.792 20.948 ;
 RECT 64.064 20.748 64.12 20.948 ;
 RECT 65.072 20.748 65.128 20.948 ;
 RECT 65.156 20.496 65.212 20.669 ;
 RECT 64.4 20.709 64.456 20.909 ;
 RECT 63.14 22.7325 63.196 22.9325 ;
 RECT 62.972 22.7325 63.028 22.9325 ;
 RECT 63.476 22.7325 63.532 22.9325 ;
 RECT 63.308 22.7325 63.364 22.9325 ;
 RECT 62.468 22.7325 62.524 22.9325 ;
 RECT 62.3 22.7325 62.356 22.9325 ;
 RECT 62.804 22.7325 62.86 22.9325 ;
 RECT 62.636 22.7325 62.692 22.9325 ;
 RECT 61.796 22.7325 61.852 22.9325 ;
 RECT 61.628 22.7325 61.684 22.9325 ;
 RECT 62.132 22.7325 62.188 22.9325 ;
 RECT 61.964 22.7325 62.02 22.9325 ;
 RECT 61.124 22.7325 61.18 22.9325 ;
 RECT 60.956 22.7325 61.012 22.9325 ;
 RECT 61.46 22.7325 61.516 22.9325 ;
 RECT 61.292 22.7325 61.348 22.9325 ;
 RECT 60.452 22.7325 60.508 22.9325 ;
 RECT 60.788 22.7325 60.844 22.9325 ;
 RECT 60.62 22.7325 60.676 22.9325 ;
 RECT 60.284 22.7325 60.34 22.9325 ;
 RECT 63.476 24.5075 63.532 24.7075 ;
 RECT 62.804 24.5075 62.86 24.7075 ;
 RECT 62.132 24.5075 62.188 24.7075 ;
 RECT 61.46 24.5075 61.516 24.7075 ;
 RECT 60.788 24.5075 60.844 24.7075 ;
 RECT 64.232 23.5045 64.288 23.7045 ;
 RECT 64.652 23.5045 64.708 23.7045 ;
 RECT 65.072 23.5045 65.128 23.7045 ;
 RECT 64.4 24.638 64.456 24.838 ;
 RECT 65.072 24.638 65.128 24.838 ;
 RECT 63.14 21.19 63.196 21.39 ;
 RECT 63.476 21.181 63.532 21.381 ;
 RECT 62.468 21.19 62.524 21.39 ;
 RECT 62.3 21.19 62.356 21.39 ;
 RECT 62.636 21.19 62.692 21.39 ;
 RECT 62.804 21.181 62.86 21.381 ;
 RECT 61.796 21.19 61.852 21.39 ;
 RECT 61.628 21.19 61.684 21.39 ;
 RECT 61.964 21.19 62.02 21.39 ;
 RECT 62.132 21.181 62.188 21.381 ;
 RECT 61.124 21.19 61.18 21.39 ;
 RECT 60.956 21.19 61.012 21.39 ;
 RECT 61.292 21.19 61.348 21.39 ;
 RECT 61.46 21.181 61.516 21.381 ;
 RECT 60.788 21.181 60.844 21.381 ;
 RECT 60.452 21.19 60.508 21.39 ;
 RECT 60.62 21.19 60.676 21.39 ;
 RECT 60.284 21.19 60.34 21.39 ;
 RECT 62.972 21.19 63.028 21.39 ;
 RECT 63.308 21.19 63.364 21.39 ;
 RECT 64.484 20.543 64.54 20.743 ;
 RECT 64.316 20.543 64.372 20.743 ;
 RECT 64.148 20.543 64.204 20.743 ;
 RECT 63.98 20.543 64.036 20.743 ;
 RECT 63.644 20.543 63.7 20.743 ;
 RECT 63.812 20.626 63.868 20.826 ;
 END
 END vss.gds2008
 PIN vss.gds2009
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.174 22.49 70.22 22.69 ;
 END
 END vss.gds2009
 PIN vss.gds2010
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.502 22.49 69.548 22.69 ;
 END
 END vss.gds2010
 PIN vss.gds2011
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.418 21.568 65.474 21.768 ;
 END
 END vss.gds2011
 PIN vss.gds2012
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.75 25.031 67.806 25.231 ;
 END
 END vss.gds2012
 PIN vss.gds2013
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.706 22.185 69.746 22.385 ;
 END
 END vss.gds2013
 PIN vss.gds2014
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.898 22.6675 69.938 22.8675 ;
 END
 END vss.gds2014
 PIN vss.gds2015
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 24.37 68.47 24.57 ;
 END
 END vss.gds2015
 PIN vss.gds2016
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 23.2245 67.302 23.4245 ;
 END
 END vss.gds2016
 PIN vss.gds2017
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.754 23.595 68.81 23.795 ;
 END
 END vss.gds2017
 PIN vss.gds2018
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 21.779 66.026 21.979 ;
 END
 END vss.gds2018
 PIN vss.gds2019
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 23.2295 68.15 23.4295 ;
 END
 END vss.gds2019
 PIN vss.gds2020
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 23.1285 66.318 23.3285 ;
 END
 END vss.gds2020
 PIN vss.gds2021
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.326 24.6335 67.382 24.8335 ;
 END
 END vss.gds2021
 PIN vss.gds2022
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 23.1945 70.086 23.3945 ;
 END
 END vss.gds2022
 PIN vss.gds2023
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 23.427 66.998 23.627 ;
 END
 END vss.gds2023
 PIN vss.gds2024
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 23.111 65.654 23.311 ;
 END
 END vss.gds2024
 PIN vss.gds2025
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 23.128 67.646 23.328 ;
 END
 END vss.gds2025
 PIN vss.gds2026
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 21.568 66.574 21.768 ;
 END
 END vss.gds2026
 PIN vss.gds2027
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 21.426 67.97 21.626 ;
 END
 END vss.gds2027
 PIN vss.gds2028
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 23.2755 68.99 23.4755 ;
 END
 END vss.gds2028
 PIN vss.gds2029
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 20.957 68.47 21.157 ;
 END
 END vss.gds2029
 PIN vss.gds2030
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 23.1945 69.414 23.3945 ;
 END
 END vss.gds2030
 PIN vss.gds2031
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 65.408 24.759 65.464 24.941 ;
 RECT 66.248 24.819 66.304 25.019 ;
 RECT 65.912 24.778 65.968 24.978 ;
 RECT 65.66 24.759 65.716 24.941 ;
 RECT 66.584 24.778 66.64 24.978 ;
 RECT 67.172 24.778 67.228 24.978 ;
 RECT 67.004 24.778 67.06 24.978 ;
 RECT 67.676 24.759 67.732 24.941 ;
 RECT 67.424 24.759 67.48 24.941 ;
 RECT 68.264 24.778 68.32 24.978 ;
 RECT 68.432 24.778 68.488 24.978 ;
 RECT 67.088 22.09 67.144 22.29 ;
 RECT 66.92 22.09 66.976 22.29 ;
 RECT 66.752 22.09 66.808 22.29 ;
 RECT 66.584 22.09 66.64 22.29 ;
 RECT 67.76 22.09 67.816 22.29 ;
 RECT 67.34 22.072 67.396 22.249 ;
 RECT 67.088 21.81 67.144 22.01 ;
 RECT 66.92 21.81 66.976 22.01 ;
 RECT 66.752 21.81 66.808 22.01 ;
 RECT 66.584 21.81 66.64 22.01 ;
 RECT 67.34 21.851 67.396 22.029 ;
 RECT 67.508 21.847 67.564 22.047 ;
 RECT 67.844 21.81 67.9 22.01 ;
 RECT 69.02 21.81 69.076 22.01 ;
 RECT 65.492 23.154 65.548 23.354 ;
 RECT 65.996 23.154 66.052 23.354 ;
 RECT 65.828 23.191 65.884 23.373 ;
 RECT 66.332 23.0835 66.388 23.2835 ;
 RECT 67.256 23.195 67.312 23.367 ;
 RECT 67.004 23.195 67.06 23.367 ;
 RECT 66.668 23.154 66.724 23.354 ;
 RECT 67.676 23.154 67.732 23.354 ;
 RECT 68.684 23.154 68.74 23.354 ;
 RECT 68.18 23.154 68.236 23.354 ;
 RECT 65.828 23.415 65.884 23.597 ;
 RECT 65.996 23.434 66.052 23.634 ;
 RECT 67.256 23.415 67.312 23.593 ;
 RECT 66.668 23.434 66.724 23.634 ;
 RECT 67.004 23.415 67.06 23.593 ;
 RECT 67.76 23.434 67.816 23.634 ;
 RECT 68.264 23.434 68.32 23.634 ;
 RECT 68.684 23.434 68.74 23.634 ;
 RECT 65.408 20.748 65.464 20.948 ;
 RECT 65.744 20.748 65.8 20.948 ;
 RECT 66.08 20.748 66.136 20.948 ;
 RECT 67.088 20.748 67.144 20.948 ;
 RECT 67.424 20.748 67.48 20.948 ;
 RECT 67.76 20.748 67.816 20.948 ;
 RECT 68.096 20.748 68.152 20.948 ;
 RECT 67.676 20.516 67.732 20.669 ;
 RECT 65.324 20.469 65.38 20.669 ;
 RECT 66.92 20.513 66.976 20.678 ;
 RECT 66.752 20.513 66.808 20.678 ;
 RECT 65.996 20.513 66.052 20.678 ;
 RECT 65.828 20.513 65.884 20.678 ;
 RECT 68.264 21.95 68.32 22.15 ;
 RECT 68.096 21.95 68.152 22.15 ;
 RECT 68.432 21.95 68.488 22.15 ;
 RECT 68.936 24.8485 68.992 25.0485 ;
 RECT 65.492 23.5045 65.548 23.7045 ;
 RECT 66.332 23.5045 66.388 23.7045 ;
 RECT 70.196 21.19 70.252 21.39 ;
 RECT 69.356 21.181 69.412 21.381 ;
 RECT 68.432 20.709 68.488 20.909 ;
 RECT 69.692 21.19 69.748 21.39 ;
 RECT 69.524 21.19 69.58 21.39 ;
 RECT 69.86 21.19 69.916 21.39 ;
 RECT 70.028 21.181 70.084 21.381 ;
 RECT 68.684 22.0615 68.74 22.2615 ;
 RECT 68.936 22.131 68.992 22.331 ;
 RECT 70.196 22.7325 70.252 22.9325 ;
 RECT 69.692 22.7325 69.748 22.9325 ;
 RECT 69.356 22.7325 69.412 22.9325 ;
 RECT 69.524 22.7325 69.58 22.9325 ;
 RECT 70.028 22.7325 70.084 22.9325 ;
 RECT 69.86 22.7325 69.916 22.9325 ;
 RECT 69.356 24.302 69.412 24.502 ;
 RECT 70.028 24.5075 70.084 24.7075 ;
 RECT 65.408 24.535 65.464 24.717 ;
 RECT 66.248 24.498 66.304 24.698 ;
 RECT 65.912 24.498 65.968 24.698 ;
 RECT 65.744 24.535 65.8 24.717 ;
 RECT 67.256 24.535 67.312 24.717 ;
 RECT 66.584 24.498 66.64 24.698 ;
 RECT 66.92 24.535 66.976 24.717 ;
 RECT 67.76 24.498 67.816 24.698 ;
 RECT 68.348 24.535 68.404 24.717 ;
 RECT 66.332 20.554 66.388 20.754 ;
 RECT 69.02 20.543 69.076 20.743 ;
 RECT 68.852 20.543 68.908 20.743 ;
 RECT 68.684 20.543 68.74 20.743 ;
 RECT 68.516 20.543 68.572 20.743 ;
 RECT 68.348 20.543 68.404 20.743 ;
 RECT 69.188 20.543 69.244 20.743 ;
 RECT 68.18 20.554 68.236 20.754 ;
 END
 END vss.gds2031
 PIN vss.gds2032
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.206 22.49 74.252 22.69 ;
 END
 END vss.gds2032
 PIN vss.gds2033
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.534 22.49 73.58 22.69 ;
 END
 END vss.gds2033
 PIN vss.gds2034
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.862 22.49 72.908 22.69 ;
 END
 END vss.gds2034
 PIN vss.gds2035
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.19 22.49 72.236 22.69 ;
 END
 END vss.gds2035
 PIN vss.gds2036
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.518 22.49 71.564 22.69 ;
 END
 END vss.gds2036
 PIN vss.gds2037
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.846 22.49 70.892 22.69 ;
 END
 END vss.gds2037
 PIN vss.gds2038
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.41 22.185 74.45 22.385 ;
 END
 END vss.gds2038
 PIN vss.gds2039
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.738 22.185 73.778 22.385 ;
 END
 END vss.gds2039
 PIN vss.gds2040
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.066 22.185 73.106 22.385 ;
 END
 END vss.gds2040
 PIN vss.gds2041
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.394 22.185 72.434 22.385 ;
 END
 END vss.gds2041
 PIN vss.gds2042
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.722 22.185 71.762 22.385 ;
 END
 END vss.gds2042
 PIN vss.gds2043
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.05 22.185 71.09 22.385 ;
 END
 END vss.gds2043
 PIN vss.gds2044
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.378 22.185 70.418 22.385 ;
 END
 END vss.gds2044
 PIN vss.gds2045
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.602 22.6675 74.642 22.8675 ;
 END
 END vss.gds2045
 PIN vss.gds2046
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.93 22.6675 73.97 22.8675 ;
 END
 END vss.gds2046
 PIN vss.gds2047
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.258 22.6675 73.298 22.8675 ;
 END
 END vss.gds2047
 PIN vss.gds2048
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.586 22.6675 72.626 22.8675 ;
 END
 END vss.gds2048
 PIN vss.gds2049
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.914 22.6675 71.954 22.8675 ;
 END
 END vss.gds2049
 PIN vss.gds2050
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.242 22.6675 71.282 22.8675 ;
 END
 END vss.gds2050
 PIN vss.gds2051
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.57 22.6675 70.61 22.8675 ;
 END
 END vss.gds2051
 PIN vss.gds2052
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 23.1945 71.43 23.3945 ;
 END
 END vss.gds2052
 PIN vss.gds2053
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 23.1945 72.102 23.3945 ;
 END
 END vss.gds2053
 PIN vss.gds2054
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 23.1945 72.774 23.3945 ;
 END
 END vss.gds2054
 PIN vss.gds2055
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 23.1945 70.758 23.3945 ;
 END
 END vss.gds2055
 PIN vss.gds2056
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 23.1945 73.446 23.3945 ;
 END
 END vss.gds2056
 PIN vss.gds2057
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 23.1945 74.118 23.3945 ;
 END
 END vss.gds2057
 PIN vss.gds2058
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 23.1945 74.79 23.3945 ;
 END
 END vss.gds2058
 PIN vss.gds2059
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 74.396 21.19 74.452 21.39 ;
 RECT 74.228 21.19 74.284 21.39 ;
 RECT 74.564 21.19 74.62 21.39 ;
 RECT 74.732 21.181 74.788 21.381 ;
 RECT 73.724 21.19 73.78 21.39 ;
 RECT 73.556 21.19 73.612 21.39 ;
 RECT 73.892 21.19 73.948 21.39 ;
 RECT 74.06 21.181 74.116 21.381 ;
 RECT 73.052 21.19 73.108 21.39 ;
 RECT 72.884 21.19 72.94 21.39 ;
 RECT 73.22 21.19 73.276 21.39 ;
 RECT 73.388 21.181 73.444 21.381 ;
 RECT 72.38 21.19 72.436 21.39 ;
 RECT 72.212 21.19 72.268 21.39 ;
 RECT 72.548 21.19 72.604 21.39 ;
 RECT 72.716 21.181 72.772 21.381 ;
 RECT 71.708 21.19 71.764 21.39 ;
 RECT 71.54 21.19 71.596 21.39 ;
 RECT 71.876 21.19 71.932 21.39 ;
 RECT 72.044 21.181 72.1 21.381 ;
 RECT 71.036 21.19 71.092 21.39 ;
 RECT 70.868 21.19 70.924 21.39 ;
 RECT 71.204 21.19 71.26 21.39 ;
 RECT 71.372 21.181 71.428 21.381 ;
 RECT 70.364 21.19 70.42 21.39 ;
 RECT 70.532 21.19 70.588 21.39 ;
 RECT 70.7 21.181 70.756 21.381 ;
 RECT 74.396 22.7325 74.452 22.9325 ;
 RECT 74.228 22.7325 74.284 22.9325 ;
 RECT 74.732 22.7325 74.788 22.9325 ;
 RECT 74.564 22.7325 74.62 22.9325 ;
 RECT 73.724 22.7325 73.78 22.9325 ;
 RECT 73.556 22.7325 73.612 22.9325 ;
 RECT 74.06 22.7325 74.116 22.9325 ;
 RECT 73.892 22.7325 73.948 22.9325 ;
 RECT 73.052 22.7325 73.108 22.9325 ;
 RECT 72.884 22.7325 72.94 22.9325 ;
 RECT 73.388 22.7325 73.444 22.9325 ;
 RECT 73.22 22.7325 73.276 22.9325 ;
 RECT 72.38 22.7325 72.436 22.9325 ;
 RECT 72.212 22.7325 72.268 22.9325 ;
 RECT 72.716 22.7325 72.772 22.9325 ;
 RECT 72.548 22.7325 72.604 22.9325 ;
 RECT 71.708 22.7325 71.764 22.9325 ;
 RECT 71.54 22.7325 71.596 22.9325 ;
 RECT 72.044 22.7325 72.1 22.9325 ;
 RECT 71.876 22.7325 71.932 22.9325 ;
 RECT 71.036 22.7325 71.092 22.9325 ;
 RECT 70.868 22.7325 70.924 22.9325 ;
 RECT 71.372 22.7325 71.428 22.9325 ;
 RECT 71.204 22.7325 71.26 22.9325 ;
 RECT 70.364 22.7325 70.42 22.9325 ;
 RECT 70.7 22.7325 70.756 22.9325 ;
 RECT 70.532 22.7325 70.588 22.9325 ;
 RECT 74.732 24.5075 74.788 24.7075 ;
 RECT 74.06 24.5075 74.116 24.7075 ;
 RECT 73.388 24.5075 73.444 24.7075 ;
 RECT 72.716 24.5075 72.772 24.7075 ;
 RECT 72.044 24.5075 72.1 24.7075 ;
 RECT 71.372 24.5075 71.428 24.7075 ;
 RECT 70.7 24.5075 70.756 24.7075 ;
 END
 END vss.gds2059
 PIN vss.gds2060
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 29.137 2.962 29.337 ;
 END
 END vss.gds2060
 PIN vss.gds2061
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 30.397 2.962 30.597 ;
 END
 END vss.gds2061
 PIN vss.gds2062
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 29.996 3.142 30.196 ;
 END
 END vss.gds2062
 PIN vss.gds2063
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.646 26.964 1.702 27.164 ;
 END
 END vss.gds2063
 PIN vss.gds2064
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.282 26.354 4.338 26.554 ;
 END
 END vss.gds2064
 PIN vss.gds2065
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 26.819 3.142 27.019 ;
 END
 END vss.gds2065
 PIN vss.gds2066
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.754 27.5075 3.794 27.7075 ;
 END
 END vss.gds2066
 PIN vss.gds2067
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 30.179 4.882 30.379 ;
 END
 END vss.gds2067
 PIN vss.gds2068
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 27.6625 5.074 27.8625 ;
 END
 END vss.gds2068
 PIN vss.gds2069
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 27.763 0.942 27.963 ;
 END
 END vss.gds2069
 PIN vss.gds2070
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 28.2545 4.194 28.4545 ;
 END
 END vss.gds2070
 PIN vss.gds2071
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 27.84 0.718 28.04 ;
 END
 END vss.gds2071
 PIN vss.gds2072
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 29.562 0.602 29.762 ;
 END
 END vss.gds2072
 PIN vss.gds2073
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 28.067 2.122 28.267 ;
 END
 END vss.gds2073
 PIN vss.gds2074
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 29.145 1.282 29.345 ;
 END
 END vss.gds2074
 PIN vss.gds2075
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 29.0745 1.462 29.2745 ;
 END
 END vss.gds2075
 PIN vss.gds2076
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 27.4095 2.302 27.6095 ;
 END
 END vss.gds2076
 PIN vss.gds2077
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 27.687 4.002 27.887 ;
 END
 END vss.gds2077
 PIN vss.gds2078
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 27.8635 5.282 28.0635 ;
 END
 END vss.gds2078
 PIN vss.gds2079
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 28.145 0.29 28.345 ;
 END
 END vss.gds2079
 PIN vss.gds2080
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 3.5 28.592 3.556 28.743 ;
 RECT 3.248 28.571 3.304 28.743 ;
 RECT 4.004 28.592 4.06 28.743 ;
 RECT 3.752 28.571 3.808 28.743 ;
 RECT 0.56 27.447 0.616 27.647 ;
 RECT 1.568 27.466 1.624 27.666 ;
 RECT 0.98 27.466 1.036 27.666 ;
 RECT 2.24 27.447 2.296 27.647 ;
 RECT 2.072 27.447 2.128 27.647 ;
 RECT 2.996 27.466 3.052 27.666 ;
 RECT 3.248 27.326 3.304 27.526 ;
 RECT 3.5 27.3245 3.556 27.5245 ;
 RECT 4.088 27.326 4.144 27.526 ;
 RECT 3.92 27.326 3.976 27.526 ;
 RECT 2.408 27.345 2.464 27.545 ;
 RECT 3.5 26.103 3.556 26.285 ;
 RECT 0.56 26.103 0.616 26.303 ;
 RECT 1.568 26.103 1.624 26.303 ;
 RECT 0.98 26.103 1.036 26.303 ;
 RECT 2.576 26.103 2.632 26.303 ;
 RECT 2.156 26.103 2.212 26.303 ;
 RECT 1.988 26.103 2.044 26.303 ;
 RECT 3.248 25.982 3.304 26.182 ;
 RECT 3.5 25.879 3.556 26.061 ;
 RECT 4.088 25.982 4.144 26.182 ;
 RECT 3.92 25.982 3.976 26.182 ;
 RECT 2.576 29.1375 2.632 29.3375 ;
 RECT 2.408 29.1375 2.464 29.3375 ;
 RECT 2.996 29.1375 3.052 29.3375 ;
 RECT 3.332 29.229 3.388 29.429 ;
 RECT 2.576 30.3975 2.632 30.5975 ;
 RECT 2.408 30.3975 2.464 30.5975 ;
 RECT 2.996 30.3975 3.052 30.5975 ;
 RECT 3.5 29.1855 3.556 29.3855 ;
 RECT 0.98 29.0525 1.036 29.2525 ;
 RECT 2.072 29.053 2.128 29.253 ;
 RECT 3.5 30.4455 3.556 30.6455 ;
 RECT 0.392 30.403 0.448 30.603 ;
 RECT 0.644 30.403 0.7 30.603 ;
 RECT 1.232 30.403 1.288 30.603 ;
 RECT 0.98 30.3125 1.036 30.5125 ;
 RECT 1.4 30.403 1.456 30.603 ;
 RECT 1.568 30.403 1.624 30.603 ;
 RECT 2.072 30.313 2.128 30.513 ;
 RECT 1.82 30.403 1.876 30.603 ;
 RECT 2.744 30.313 2.8 30.513 ;
 RECT 3.164 30.403 3.22 30.603 ;
 RECT 2.24 30.403 2.296 30.603 ;
 RECT 0.392 29.143 0.448 29.343 ;
 RECT 0.812 29.229 0.868 29.429 ;
 RECT 0.644 29.143 0.7 29.343 ;
 RECT 1.232 29.143 1.288 29.343 ;
 RECT 1.4 29.143 1.456 29.343 ;
 RECT 1.568 29.143 1.624 29.343 ;
 RECT 1.82 29.143 1.876 29.343 ;
 RECT 2.24 29.143 2.296 29.343 ;
 RECT 2.744 29.053 2.8 29.253 ;
 RECT 3.164 29.143 3.22 29.343 ;
 RECT 3.92 30.403 3.976 30.603 ;
 RECT 3.92 29.143 3.976 29.343 ;
 RECT 3.752 29.413 3.808 29.613 ;
 RECT 4.508 29.3425 4.564 29.5425 ;
 RECT 0.56 25.7715 0.616 25.9715 ;
 RECT 1.568 25.7715 1.624 25.9715 ;
 RECT 0.98 25.7715 1.036 25.9715 ;
 RECT 2.072 25.842 2.128 26.042 ;
 RECT 1.904 25.842 1.96 26.042 ;
 RECT 3.08 25.842 3.136 26.042 ;
 RECT 2.912 25.842 2.968 26.042 ;
 RECT 2.744 25.842 2.8 26.042 ;
 RECT 4.676 25.982 4.732 26.182 ;
 RECT 4.424 25.9765 4.48 26.1765 ;
 RECT 1.568 27.1155 1.624 27.3155 ;
 RECT 0.98 27.1155 1.036 27.3155 ;
 RECT 0.56 27.166 0.616 27.366 ;
 RECT 2.156 27.205 2.212 27.405 ;
 RECT 1.988 27.186 2.044 27.386 ;
 RECT 2.996 27.186 3.052 27.386 ;
 RECT 4.676 27.326 4.732 27.526 ;
 RECT 4.424 27.326 4.48 27.526 ;
 RECT 2.744 27.326 2.8 27.526 ;
 RECT 0.56 28.549 0.616 28.749 ;
 RECT 1.568 28.549 1.624 28.749 ;
 RECT 0.98 28.549 1.036 28.749 ;
 RECT 1.988 28.528 2.044 28.728 ;
 RECT 2.492 28.528 2.548 28.728 ;
 RECT 2.24 28.528 2.296 28.728 ;
 RECT 2.744 28.528 2.8 28.728 ;
 RECT 2.996 28.528 3.052 28.728 ;
 RECT 4.676 28.528 4.732 28.728 ;
 RECT 4.424 28.528 4.48 28.728 ;
 END
 END vss.gds2080
 PIN vss.gds2081
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.046 25.982 10.086 26.182 ;
 END
 END vss.gds2081
 PIN vss.gds2082
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.374 25.982 9.414 26.182 ;
 END
 END vss.gds2082
 PIN vss.gds2083
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.702 25.982 8.742 26.182 ;
 END
 END vss.gds2083
 PIN vss.gds2084
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.03 25.982 8.07 26.182 ;
 END
 END vss.gds2084
 PIN vss.gds2085
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.778 25.775 9.824 25.975 ;
 END
 END vss.gds2085
 PIN vss.gds2086
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.174 25.775 10.214 25.975 ;
 END
 END vss.gds2086
 PIN vss.gds2087
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.106 25.775 9.152 25.975 ;
 END
 END vss.gds2087
 PIN vss.gds2088
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.502 25.775 9.542 25.975 ;
 END
 END vss.gds2088
 PIN vss.gds2089
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.434 25.775 8.48 25.975 ;
 END
 END vss.gds2089
 PIN vss.gds2090
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.83 25.775 8.87 25.975 ;
 END
 END vss.gds2090
 PIN vss.gds2091
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.762 25.775 7.808 25.975 ;
 END
 END vss.gds2091
 PIN vss.gds2092
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.158 25.775 8.198 25.975 ;
 END
 END vss.gds2092
 PIN vss.gds2093
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.09 25.775 7.136 25.975 ;
 END
 END vss.gds2093
 PIN vss.gds2094
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.486 25.775 7.526 25.975 ;
 END
 END vss.gds2094
 PIN vss.gds2095
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.358 25.982 7.398 26.182 ;
 END
 END vss.gds2095
 PIN vss.gds2096
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 28.2535 9.69 28.4535 ;
 END
 END vss.gds2096
 PIN vss.gds2097
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 28.2535 9.018 28.4535 ;
 END
 END vss.gds2097
 PIN vss.gds2098
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.942 26.9135 7.002 27.1135 ;
 END
 END vss.gds2098
 PIN vss.gds2099
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.734 26.9905 6.774 27.1905 ;
 END
 END vss.gds2099
 PIN vss.gds2100
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.606 26.9905 6.646 27.1905 ;
 END
 END vss.gds2100
 PIN vss.gds2101
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 28.079 6.178 28.279 ;
 END
 END vss.gds2101
 PIN vss.gds2102
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 27.6625 5.474 27.8625 ;
 END
 END vss.gds2102
 PIN vss.gds2103
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 28.2535 8.346 28.4535 ;
 END
 END vss.gds2103
 PIN vss.gds2104
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 28.2535 7.674 28.4535 ;
 END
 END vss.gds2104
 PIN vss.gds2105
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 27.7585 5.73 27.9585 ;
 END
 END vss.gds2105
 PIN vss.gds2106
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 27.6625 5.986 27.8625 ;
 END
 END vss.gds2106
 PIN vss.gds2107
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 28.326 6.434 28.526 ;
 END
 END vss.gds2107
 PIN vss.gds2108
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 10.136 28.573 10.192 28.773 ;
 RECT 9.632 28.563 9.688 28.763 ;
 RECT 9.464 28.573 9.52 28.773 ;
 RECT 8.96 28.563 9.016 28.763 ;
 RECT 8.792 28.573 8.848 28.773 ;
 RECT 8.288 28.563 8.344 28.763 ;
 RECT 8.12 28.573 8.176 28.773 ;
 RECT 6.944 28.563 7 28.763 ;
 RECT 7.616 28.563 7.672 28.763 ;
 RECT 7.448 28.573 7.504 28.773 ;
 RECT 5.6 27.466 5.656 27.666 ;
 RECT 9.968 25.801 10.024 26.001 ;
 RECT 9.8 25.801 9.856 26.001 ;
 RECT 10.136 25.816 10.192 26.016 ;
 RECT 9.296 25.801 9.352 26.001 ;
 RECT 9.128 25.801 9.184 26.001 ;
 RECT 9.464 25.816 9.52 26.016 ;
 RECT 9.632 25.816 9.688 26.016 ;
 RECT 8.624 25.801 8.68 26.001 ;
 RECT 8.456 25.801 8.512 26.001 ;
 RECT 8.792 25.816 8.848 26.016 ;
 RECT 8.96 25.816 9.016 26.016 ;
 RECT 7.952 25.801 8.008 26.001 ;
 RECT 7.784 25.801 7.84 26.001 ;
 RECT 8.12 25.816 8.176 26.016 ;
 RECT 8.288 25.816 8.344 26.016 ;
 RECT 7.28 25.801 7.336 26.001 ;
 RECT 7.112 25.801 7.168 26.001 ;
 RECT 6.944 25.816 7 26.016 ;
 RECT 7.448 25.816 7.504 26.016 ;
 RECT 7.616 25.816 7.672 26.016 ;
 RECT 9.968 26.875 10.024 27.075 ;
 RECT 9.8 26.875 9.856 27.075 ;
 RECT 10.136 26.875 10.192 27.075 ;
 RECT 9.296 26.875 9.352 27.075 ;
 RECT 9.128 26.875 9.184 27.075 ;
 RECT 9.632 26.875 9.688 27.075 ;
 RECT 9.464 26.875 9.52 27.075 ;
 RECT 8.624 26.875 8.68 27.075 ;
 RECT 8.456 26.875 8.512 27.075 ;
 RECT 8.96 26.875 9.016 27.075 ;
 RECT 8.792 26.875 8.848 27.075 ;
 RECT 7.952 26.875 8.008 27.075 ;
 RECT 7.784 26.875 7.84 27.075 ;
 RECT 8.288 26.875 8.344 27.075 ;
 RECT 8.12 26.875 8.176 27.075 ;
 RECT 7.28 26.875 7.336 27.075 ;
 RECT 6.944 26.875 7 27.075 ;
 RECT 7.112 26.875 7.168 27.075 ;
 RECT 7.616 26.875 7.672 27.075 ;
 RECT 7.448 26.875 7.504 27.075 ;
 RECT 6.524 30.396 6.58 30.596 ;
 RECT 6.692 29.286 6.748 29.486 ;
 RECT 6.524 29.136 6.58 29.336 ;
 RECT 6.608 29.413 6.664 29.613 ;
 RECT 5.432 25.982 5.488 26.182 ;
 RECT 5.6 25.982 5.656 26.182 ;
 RECT 5.768 25.982 5.824 26.182 ;
 RECT 5.936 25.982 5.992 26.182 ;
 RECT 6.44 25.982 6.496 26.182 ;
 RECT 6.104 25.982 6.16 26.182 ;
 RECT 6.272 25.982 6.328 26.182 ;
 RECT 5.432 27.326 5.488 27.526 ;
 RECT 5.6 27.186 5.656 27.386 ;
 RECT 5.768 27.326 5.824 27.526 ;
 RECT 5.936 27.326 5.992 27.526 ;
 RECT 6.104 27.326 6.16 27.526 ;
 RECT 6.272 27.326 6.328 27.526 ;
 RECT 6.44 27.326 6.496 27.526 ;
 RECT 5.432 28.528 5.488 28.728 ;
 RECT 5.6 28.528 5.656 28.728 ;
 RECT 5.768 28.528 5.824 28.728 ;
 RECT 5.936 28.528 5.992 28.728 ;
 RECT 6.104 28.528 6.16 28.728 ;
 RECT 6.272 28.528 6.328 28.728 ;
 RECT 6.44 28.528 6.496 28.728 ;
 END
 END vss.gds2108
 PIN vss.gds2109
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.262 26.9905 14.318 27.1905 ;
 END
 END vss.gds2109
 PIN vss.gds2110
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 29.682 14.87 29.882 ;
 END
 END vss.gds2110
 PIN vss.gds2111
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 26.4595 13.898 26.6595 ;
 END
 END vss.gds2111
 PIN vss.gds2112
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.062 25.982 12.102 26.182 ;
 END
 END vss.gds2112
 PIN vss.gds2113
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.39 25.982 11.43 26.182 ;
 END
 END vss.gds2113
 PIN vss.gds2114
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.718 25.982 10.758 26.182 ;
 END
 END vss.gds2114
 PIN vss.gds2115
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 26.2765 14.87 26.4765 ;
 END
 END vss.gds2115
 PIN vss.gds2116
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 26.102 13.058 26.302 ;
 END
 END vss.gds2116
 PIN vss.gds2117
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.794 25.775 11.84 25.975 ;
 END
 END vss.gds2117
 PIN vss.gds2118
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.19 25.775 12.23 25.975 ;
 END
 END vss.gds2118
 PIN vss.gds2119
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.122 25.775 11.168 25.975 ;
 END
 END vss.gds2119
 PIN vss.gds2120
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.518 25.775 11.558 25.975 ;
 END
 END vss.gds2120
 PIN vss.gds2121
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.45 25.775 10.496 25.975 ;
 END
 END vss.gds2121
 PIN vss.gds2122
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.846 25.775 10.886 25.975 ;
 END
 END vss.gds2122
 PIN vss.gds2123
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.262 29.231 13.318 29.431 ;
 END
 END vss.gds2123
 PIN vss.gds2124
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 28.2535 11.706 28.4535 ;
 END
 END vss.gds2124
 PIN vss.gds2125
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 28.2535 11.034 28.4535 ;
 END
 END vss.gds2125
 PIN vss.gds2126
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 28.2535 10.362 28.4535 ;
 END
 END vss.gds2126
 PIN vss.gds2127
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 28.4415 15.162 28.6415 ;
 END
 END vss.gds2127
 PIN vss.gds2128
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 29.642 13.898 29.842 ;
 END
 END vss.gds2128
 PIN vss.gds2129
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 28.5025 14.498 28.7025 ;
 END
 END vss.gds2129
 PIN vss.gds2130
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 28.2885 13.658 28.4885 ;
 END
 END vss.gds2130
 PIN vss.gds2131
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 27.837 12.378 28.037 ;
 END
 END vss.gds2131
 PIN vss.gds2132
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 27.6625 12.59 27.8625 ;
 END
 END vss.gds2132
 PIN vss.gds2133
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 28.3975 12.818 28.5975 ;
 END
 END vss.gds2133
 PIN vss.gds2134
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 13.244 28.469 13.3 28.669 ;
 RECT 12.32 28.563 12.376 28.763 ;
 RECT 12.152 28.573 12.208 28.773 ;
 RECT 11.648 28.563 11.704 28.763 ;
 RECT 11.48 28.573 11.536 28.773 ;
 RECT 10.976 28.563 11.032 28.763 ;
 RECT 10.808 28.573 10.864 28.773 ;
 RECT 10.304 28.563 10.36 28.763 ;
 RECT 12.824 26.122 12.88 26.322 ;
 RECT 15.176 26.122 15.232 26.322 ;
 RECT 15.008 26.122 15.064 26.322 ;
 RECT 13.664 26.103 13.72 26.303 ;
 RECT 12.992 26.103 13.048 26.303 ;
 RECT 13.16 26.103 13.216 26.303 ;
 RECT 13.496 26.103 13.552 26.303 ;
 RECT 14 26.103 14.056 26.303 ;
 RECT 14.168 26.103 14.224 26.303 ;
 RECT 13.832 26.103 13.888 26.303 ;
 RECT 14.84 26.103 14.896 26.303 ;
 RECT 14.504 26.122 14.56 26.322 ;
 RECT 14.672 26.122 14.728 26.322 ;
 RECT 13.244 25.842 13.3 26.042 ;
 RECT 13.58 25.842 13.636 26.042 ;
 RECT 12.908 25.842 12.964 26.042 ;
 RECT 13.916 25.842 13.972 26.042 ;
 RECT 14.252 25.842 14.308 26.042 ;
 RECT 14.924 25.842 14.98 26.042 ;
 RECT 11.984 25.801 12.04 26.001 ;
 RECT 11.816 25.801 11.872 26.001 ;
 RECT 12.152 25.816 12.208 26.016 ;
 RECT 12.32 25.816 12.376 26.016 ;
 RECT 11.312 25.801 11.368 26.001 ;
 RECT 11.144 25.801 11.2 26.001 ;
 RECT 11.48 25.816 11.536 26.016 ;
 RECT 11.648 25.816 11.704 26.016 ;
 RECT 10.64 25.801 10.696 26.001 ;
 RECT 10.472 25.801 10.528 26.001 ;
 RECT 10.808 25.816 10.864 26.016 ;
 RECT 10.976 25.816 11.032 26.016 ;
 RECT 10.304 25.816 10.36 26.016 ;
 RECT 14 29.82 14.056 29.993 ;
 RECT 14.168 29.793 14.224 29.993 ;
 RECT 14.336 30.413 14.392 30.613 ;
 RECT 14.168 30.413 14.224 30.613 ;
 RECT 13.16 27.459 13.216 27.659 ;
 RECT 13.412 27.673 13.468 27.873 ;
 RECT 14.336 29.153 14.392 29.353 ;
 RECT 14.168 29.153 14.224 29.353 ;
 RECT 15.008 29.363 15.064 29.563 ;
 RECT 14.84 29.837 14.896 30.002 ;
 RECT 14.672 29.837 14.728 30.002 ;
 RECT 11.984 26.875 12.04 27.075 ;
 RECT 11.816 26.875 11.872 27.075 ;
 RECT 12.32 26.875 12.376 27.075 ;
 RECT 12.152 26.875 12.208 27.075 ;
 RECT 11.312 26.875 11.368 27.075 ;
 RECT 11.144 26.875 11.2 27.075 ;
 RECT 11.648 26.875 11.704 27.075 ;
 RECT 11.48 26.875 11.536 27.075 ;
 RECT 10.64 26.875 10.696 27.075 ;
 RECT 10.472 26.875 10.528 27.075 ;
 RECT 10.976 26.875 11.032 27.075 ;
 RECT 10.808 26.875 10.864 27.075 ;
 RECT 10.304 26.875 10.36 27.075 ;
 RECT 13.664 29.287 13.72 29.487 ;
 END
 END vss.gds2134
 PIN vss.gds2135
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.958 25.982 19.998 26.182 ;
 END
 END vss.gds2135
 PIN vss.gds2136
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.286 25.982 19.326 26.182 ;
 END
 END vss.gds2136
 PIN vss.gds2137
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.614 25.982 18.654 26.182 ;
 END
 END vss.gds2137
 PIN vss.gds2138
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.69 25.775 19.736 25.975 ;
 END
 END vss.gds2138
 PIN vss.gds2139
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.086 25.775 20.126 25.975 ;
 END
 END vss.gds2139
 PIN vss.gds2140
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 26.2765 16.146 26.4765 ;
 END
 END vss.gds2140
 PIN vss.gds2141
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 30.197 15.418 30.397 ;
 END
 END vss.gds2141
 PIN vss.gds2142
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.438 29.023 17.494 29.223 ;
 END
 END vss.gds2142
 PIN vss.gds2143
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 28.2535 20.274 28.4535 ;
 END
 END vss.gds2143
 PIN vss.gds2144
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.018 25.775 19.064 25.975 ;
 END
 END vss.gds2144
 PIN vss.gds2145
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.414 25.775 19.454 25.975 ;
 END
 END vss.gds2145
 PIN vss.gds2146
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.346 25.775 18.392 25.975 ;
 END
 END vss.gds2146
 PIN vss.gds2147
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.742 25.775 18.782 25.975 ;
 END
 END vss.gds2147
 PIN vss.gds2148
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 26.52 16.814 26.72 ;
 END
 END vss.gds2148
 PIN vss.gds2149
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 30.397 16.146 30.597 ;
 END
 END vss.gds2149
 PIN vss.gds2150
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 29.137 16.146 29.337 ;
 END
 END vss.gds2150
 PIN vss.gds2151
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 30.0685 17.314 30.2685 ;
 END
 END vss.gds2151
 PIN vss.gds2152
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 28.2535 18.93 28.4535 ;
 END
 END vss.gds2152
 PIN vss.gds2153
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 28.2535 19.602 28.4535 ;
 END
 END vss.gds2153
 PIN vss.gds2154
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 28.224 16.994 28.424 ;
 END
 END vss.gds2154
 PIN vss.gds2155
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 28.5025 15.842 28.7025 ;
 END
 END vss.gds2155
 PIN vss.gds2156
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 27.837 18.258 28.037 ;
 END
 END vss.gds2156
 PIN vss.gds2157
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 28.3975 17.834 28.5975 ;
 END
 END vss.gds2157
 PIN vss.gds2158
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 28.277 16.49 28.477 ;
 END
 END vss.gds2158
 PIN vss.gds2159
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 20.216 28.563 20.272 28.763 ;
 RECT 20.048 28.573 20.104 28.773 ;
 RECT 19.544 28.563 19.6 28.763 ;
 RECT 19.376 28.573 19.432 28.773 ;
 RECT 18.2 28.563 18.256 28.763 ;
 RECT 18.872 28.563 18.928 28.763 ;
 RECT 18.704 28.573 18.76 28.773 ;
 RECT 16.1 26.122 16.156 26.322 ;
 RECT 15.596 26.122 15.652 26.322 ;
 RECT 15.428 26.122 15.484 26.322 ;
 RECT 15.764 26.122 15.82 26.322 ;
 RECT 16.604 26.122 16.66 26.322 ;
 RECT 16.772 26.122 16.828 26.322 ;
 RECT 16.436 26.122 16.492 26.322 ;
 RECT 16.268 26.122 16.324 26.322 ;
 RECT 17.696 26.122 17.752 26.322 ;
 RECT 17.276 26.103 17.332 26.285 ;
 RECT 17.024 26.103 17.08 26.285 ;
 RECT 19.88 25.801 19.936 26.001 ;
 RECT 19.712 25.801 19.768 26.001 ;
 RECT 20.048 25.816 20.104 26.016 ;
 RECT 20.216 25.816 20.272 26.016 ;
 RECT 15.26 25.842 15.316 26.042 ;
 RECT 15.596 25.842 15.652 26.042 ;
 RECT 15.932 25.842 15.988 26.042 ;
 RECT 16.268 25.842 16.324 26.042 ;
 RECT 17.192 25.879 17.248 26.061 ;
 RECT 16.94 25.879 16.996 26.061 ;
 RECT 17.528 25.842 17.584 26.042 ;
 RECT 17.78 25.842 17.836 26.042 ;
 RECT 19.208 25.801 19.264 26.001 ;
 RECT 19.04 25.801 19.096 26.001 ;
 RECT 19.376 25.816 19.432 26.016 ;
 RECT 19.544 25.816 19.6 26.016 ;
 RECT 18.2 25.816 18.256 26.016 ;
 RECT 18.704 25.816 18.76 26.016 ;
 RECT 18.872 25.816 18.928 26.016 ;
 RECT 15.596 28.804 15.652 29.004 ;
 RECT 15.848 28.807 15.904 29.007 ;
 RECT 16.52 29.84 16.576 29.993 ;
 RECT 15.764 29.837 15.82 30.002 ;
 RECT 15.596 29.837 15.652 30.002 ;
 RECT 15.596 30.064 15.652 30.264 ;
 RECT 15.848 30.067 15.904 30.267 ;
 RECT 18.536 25.801 18.592 26.001 ;
 RECT 18.368 25.801 18.424 26.001 ;
 RECT 18.116 26.654 18.172 26.854 ;
 RECT 15.428 29.363 15.484 29.563 ;
 RECT 16.856 29.2115 16.912 29.4115 ;
 RECT 16.352 29.4635 16.408 29.6635 ;
 RECT 19.88 26.875 19.936 27.075 ;
 RECT 19.712 26.875 19.768 27.075 ;
 RECT 20.216 26.875 20.272 27.075 ;
 RECT 20.048 26.875 20.104 27.075 ;
 RECT 19.208 26.875 19.264 27.075 ;
 RECT 19.04 26.875 19.096 27.075 ;
 RECT 19.544 26.875 19.6 27.075 ;
 RECT 19.376 26.875 19.432 27.075 ;
 RECT 18.536 26.875 18.592 27.075 ;
 RECT 18.2 26.875 18.256 27.075 ;
 RECT 18.368 26.875 18.424 27.075 ;
 RECT 18.872 26.875 18.928 27.075 ;
 RECT 18.704 26.875 18.76 27.075 ;
 END
 END vss.gds2159
 PIN vss.gds2160
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.082 25.982 25.122 26.182 ;
 END
 END vss.gds2160
 PIN vss.gds2161
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.41 25.982 24.45 26.182 ;
 END
 END vss.gds2161
 PIN vss.gds2162
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.318 25.982 23.358 26.182 ;
 END
 END vss.gds2162
 PIN vss.gds2163
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.646 25.982 22.686 26.182 ;
 END
 END vss.gds2163
 PIN vss.gds2164
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.974 25.982 22.014 26.182 ;
 END
 END vss.gds2164
 PIN vss.gds2165
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.302 25.982 21.342 26.182 ;
 END
 END vss.gds2165
 PIN vss.gds2166
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.63 25.982 20.67 26.182 ;
 END
 END vss.gds2166
 PIN vss.gds2167
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.814 25.775 24.86 25.975 ;
 END
 END vss.gds2167
 PIN vss.gds2168
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.21 25.775 25.25 25.975 ;
 END
 END vss.gds2168
 PIN vss.gds2169
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.142 25.775 24.188 25.975 ;
 END
 END vss.gds2169
 PIN vss.gds2170
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.538 25.775 24.578 25.975 ;
 END
 END vss.gds2170
 PIN vss.gds2171
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.05 25.775 23.096 25.975 ;
 END
 END vss.gds2171
 PIN vss.gds2172
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.446 25.775 23.486 25.975 ;
 END
 END vss.gds2172
 PIN vss.gds2173
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.378 25.775 22.424 25.975 ;
 END
 END vss.gds2173
 PIN vss.gds2174
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.774 25.775 22.814 25.975 ;
 END
 END vss.gds2174
 PIN vss.gds2175
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.706 25.775 21.752 25.975 ;
 END
 END vss.gds2175
 PIN vss.gds2176
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.102 25.775 22.142 25.975 ;
 END
 END vss.gds2176
 PIN vss.gds2177
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.034 25.775 21.08 25.975 ;
 END
 END vss.gds2177
 PIN vss.gds2178
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.43 25.775 21.47 25.975 ;
 END
 END vss.gds2178
 PIN vss.gds2179
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.362 25.775 20.408 25.975 ;
 END
 END vss.gds2179
 PIN vss.gds2180
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.758 25.775 20.798 25.975 ;
 END
 END vss.gds2180
 PIN vss.gds2181
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.722 26.9905 23.762 27.1905 ;
 END
 END vss.gds2181
 PIN vss.gds2182
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.866 26.9905 23.906 27.1905 ;
 END
 END vss.gds2182
 PIN vss.gds2183
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 28.2535 24.726 28.4535 ;
 END
 END vss.gds2183
 PIN vss.gds2184
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 28.2535 21.618 28.4535 ;
 END
 END vss.gds2184
 PIN vss.gds2185
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.994 26.9135 24.054 27.1135 ;
 END
 END vss.gds2185
 PIN vss.gds2186
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 28.2535 20.946 28.4535 ;
 END
 END vss.gds2186
 PIN vss.gds2187
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 28.2535 22.29 28.4535 ;
 END
 END vss.gds2187
 PIN vss.gds2188
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 28.2535 22.962 28.4535 ;
 END
 END vss.gds2188
 PIN vss.gds2189
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 28.2535 23.634 28.4535 ;
 END
 END vss.gds2189
 PIN vss.gds2190
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 25.172 28.573 25.228 28.773 ;
 RECT 23.996 28.563 24.052 28.763 ;
 RECT 24.668 28.563 24.724 28.763 ;
 RECT 24.5 28.573 24.556 28.773 ;
 RECT 23.576 28.563 23.632 28.763 ;
 RECT 23.408 28.573 23.464 28.773 ;
 RECT 22.904 28.563 22.96 28.763 ;
 RECT 22.736 28.573 22.792 28.773 ;
 RECT 22.232 28.563 22.288 28.763 ;
 RECT 22.064 28.573 22.12 28.773 ;
 RECT 21.56 28.563 21.616 28.763 ;
 RECT 21.392 28.573 21.448 28.773 ;
 RECT 20.888 28.563 20.944 28.763 ;
 RECT 20.72 28.573 20.776 28.773 ;
 RECT 25.004 25.801 25.06 26.001 ;
 RECT 24.836 25.801 24.892 26.001 ;
 RECT 25.172 25.816 25.228 26.016 ;
 RECT 23.996 25.816 24.052 26.016 ;
 RECT 24.5 25.816 24.556 26.016 ;
 RECT 24.668 25.816 24.724 26.016 ;
 RECT 23.408 25.816 23.464 26.016 ;
 RECT 23.576 25.816 23.632 26.016 ;
 RECT 22.568 25.801 22.624 26.001 ;
 RECT 22.4 25.801 22.456 26.001 ;
 RECT 22.736 25.816 22.792 26.016 ;
 RECT 22.904 25.816 22.96 26.016 ;
 RECT 21.896 25.801 21.952 26.001 ;
 RECT 21.728 25.801 21.784 26.001 ;
 RECT 22.064 25.816 22.12 26.016 ;
 RECT 22.232 25.816 22.288 26.016 ;
 RECT 21.224 25.801 21.28 26.001 ;
 RECT 21.056 25.801 21.112 26.001 ;
 RECT 21.392 25.816 21.448 26.016 ;
 RECT 21.56 25.816 21.616 26.016 ;
 RECT 20.72 25.816 20.776 26.016 ;
 RECT 20.888 25.816 20.944 26.016 ;
 RECT 20.552 25.801 20.608 26.001 ;
 RECT 20.384 25.801 20.44 26.001 ;
 RECT 24.332 25.801 24.388 26.001 ;
 RECT 24.164 25.801 24.22 26.001 ;
 RECT 23.24 25.801 23.296 26.001 ;
 RECT 23.072 25.801 23.128 26.001 ;
 RECT 23.912 29.3 23.968 29.5 ;
 RECT 25.004 26.875 25.06 27.075 ;
 RECT 24.836 26.875 24.892 27.075 ;
 RECT 25.172 26.875 25.228 27.075 ;
 RECT 24.332 26.875 24.388 27.075 ;
 RECT 23.996 26.875 24.052 27.075 ;
 RECT 24.164 26.875 24.22 27.075 ;
 RECT 24.668 26.875 24.724 27.075 ;
 RECT 24.5 26.875 24.556 27.075 ;
 RECT 23.24 26.875 23.296 27.075 ;
 RECT 23.072 26.875 23.128 27.075 ;
 RECT 23.576 26.875 23.632 27.075 ;
 RECT 23.408 26.875 23.464 27.075 ;
 RECT 22.568 26.875 22.624 27.075 ;
 RECT 22.4 26.875 22.456 27.075 ;
 RECT 22.904 26.875 22.96 27.075 ;
 RECT 22.736 26.875 22.792 27.075 ;
 RECT 21.896 26.875 21.952 27.075 ;
 RECT 21.728 26.875 21.784 27.075 ;
 RECT 22.232 26.875 22.288 27.075 ;
 RECT 22.064 26.875 22.12 27.075 ;
 RECT 21.224 26.875 21.28 27.075 ;
 RECT 21.056 26.875 21.112 27.075 ;
 RECT 21.56 26.875 21.616 27.075 ;
 RECT 21.392 26.875 21.448 27.075 ;
 RECT 20.552 26.875 20.608 27.075 ;
 RECT 20.888 26.875 20.944 27.075 ;
 RECT 20.72 26.875 20.776 27.075 ;
 RECT 20.384 26.875 20.44 27.075 ;
 RECT 23.744 28.7285 23.8 28.9285 ;
 END
 END vss.gds2190
 PIN vss.gds2191
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.114 25.982 29.154 26.182 ;
 END
 END vss.gds2191
 PIN vss.gds2192
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.442 25.982 28.482 26.182 ;
 END
 END vss.gds2192
 PIN vss.gds2193
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.77 25.982 27.81 26.182 ;
 END
 END vss.gds2193
 PIN vss.gds2194
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.098 25.982 27.138 26.182 ;
 END
 END vss.gds2194
 PIN vss.gds2195
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.426 25.982 26.466 26.182 ;
 END
 END vss.gds2195
 PIN vss.gds2196
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.754 25.982 25.794 26.182 ;
 END
 END vss.gds2196
 PIN vss.gds2197
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.846 25.775 28.892 25.975 ;
 END
 END vss.gds2197
 PIN vss.gds2198
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.242 25.775 29.282 25.975 ;
 END
 END vss.gds2198
 PIN vss.gds2199
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.174 25.775 28.22 25.975 ;
 END
 END vss.gds2199
 PIN vss.gds2200
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.57 25.775 28.61 25.975 ;
 END
 END vss.gds2200
 PIN vss.gds2201
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.502 25.775 27.548 25.975 ;
 END
 END vss.gds2201
 PIN vss.gds2202
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.898 25.775 27.938 25.975 ;
 END
 END vss.gds2202
 PIN vss.gds2203
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.83 25.775 26.876 25.975 ;
 END
 END vss.gds2203
 PIN vss.gds2204
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.226 25.775 27.266 25.975 ;
 END
 END vss.gds2204
 PIN vss.gds2205
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.158 25.775 26.204 25.975 ;
 END
 END vss.gds2205
 PIN vss.gds2206
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.554 25.775 26.594 25.975 ;
 END
 END vss.gds2206
 PIN vss.gds2207
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.486 25.775 25.532 25.975 ;
 END
 END vss.gds2207
 PIN vss.gds2208
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.882 25.775 25.922 25.975 ;
 END
 END vss.gds2208
 PIN vss.gds2209
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 28.2535 28.758 28.4535 ;
 END
 END vss.gds2209
 PIN vss.gds2210
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 28.2535 28.086 28.4535 ;
 END
 END vss.gds2210
 PIN vss.gds2211
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 28.2535 27.414 28.4535 ;
 END
 END vss.gds2211
 PIN vss.gds2212
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 28.2535 26.742 28.4535 ;
 END
 END vss.gds2212
 PIN vss.gds2213
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 28.2535 26.07 28.4535 ;
 END
 END vss.gds2213
 PIN vss.gds2214
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 28.2535 25.398 28.4535 ;
 END
 END vss.gds2214
 PIN vss.gds2215
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 27.837 29.43 28.037 ;
 END
 END vss.gds2215
 PIN vss.gds2216
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 26.102 30.11 26.302 ;
 END
 END vss.gds2216
 PIN vss.gds2217
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 28.3975 29.87 28.5975 ;
 END
 END vss.gds2217
 PIN vss.gds2218
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 27.6625 29.642 27.8625 ;
 END
 END vss.gds2218
 PIN vss.gds2219
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.372 28.563 29.428 28.763 ;
 RECT 29.204 28.573 29.26 28.773 ;
 RECT 28.7 28.563 28.756 28.763 ;
 RECT 28.532 28.573 28.588 28.773 ;
 RECT 28.028 28.563 28.084 28.763 ;
 RECT 27.86 28.573 27.916 28.773 ;
 RECT 27.356 28.563 27.412 28.763 ;
 RECT 27.188 28.573 27.244 28.773 ;
 RECT 26.684 28.563 26.74 28.763 ;
 RECT 26.516 28.573 26.572 28.773 ;
 RECT 26.012 28.563 26.068 28.763 ;
 RECT 25.844 28.573 25.9 28.773 ;
 RECT 25.34 28.563 25.396 28.763 ;
 RECT 29.876 26.122 29.932 26.322 ;
 RECT 30.044 26.103 30.1 26.303 ;
 RECT 30.212 26.103 30.268 26.303 ;
 RECT 29.96 25.842 30.016 26.042 ;
 RECT 29.036 25.801 29.092 26.001 ;
 RECT 28.868 25.801 28.924 26.001 ;
 RECT 29.204 25.816 29.26 26.016 ;
 RECT 29.372 25.816 29.428 26.016 ;
 RECT 28.364 25.801 28.42 26.001 ;
 RECT 28.196 25.801 28.252 26.001 ;
 RECT 28.532 25.816 28.588 26.016 ;
 RECT 28.7 25.816 28.756 26.016 ;
 RECT 27.692 25.801 27.748 26.001 ;
 RECT 27.524 25.801 27.58 26.001 ;
 RECT 27.86 25.816 27.916 26.016 ;
 RECT 28.028 25.816 28.084 26.016 ;
 RECT 27.02 25.801 27.076 26.001 ;
 RECT 26.852 25.801 26.908 26.001 ;
 RECT 27.188 25.816 27.244 26.016 ;
 RECT 27.356 25.816 27.412 26.016 ;
 RECT 26.348 25.801 26.404 26.001 ;
 RECT 26.18 25.801 26.236 26.001 ;
 RECT 26.516 25.816 26.572 26.016 ;
 RECT 26.684 25.816 26.74 26.016 ;
 RECT 25.676 25.801 25.732 26.001 ;
 RECT 25.508 25.801 25.564 26.001 ;
 RECT 25.844 25.816 25.9 26.016 ;
 RECT 26.012 25.816 26.068 26.016 ;
 RECT 25.34 25.816 25.396 26.016 ;
 RECT 30.212 27.459 30.268 27.659 ;
 RECT 29.036 26.875 29.092 27.075 ;
 RECT 28.868 26.875 28.924 27.075 ;
 RECT 29.372 26.875 29.428 27.075 ;
 RECT 29.204 26.875 29.26 27.075 ;
 RECT 28.364 26.875 28.42 27.075 ;
 RECT 28.196 26.875 28.252 27.075 ;
 RECT 28.7 26.875 28.756 27.075 ;
 RECT 28.532 26.875 28.588 27.075 ;
 RECT 27.692 26.875 27.748 27.075 ;
 RECT 27.524 26.875 27.58 27.075 ;
 RECT 28.028 26.875 28.084 27.075 ;
 RECT 27.86 26.875 27.916 27.075 ;
 RECT 27.02 26.875 27.076 27.075 ;
 RECT 26.852 26.875 26.908 27.075 ;
 RECT 27.356 26.875 27.412 27.075 ;
 RECT 27.188 26.875 27.244 27.075 ;
 RECT 26.348 26.875 26.404 27.075 ;
 RECT 26.18 26.875 26.236 27.075 ;
 RECT 26.684 26.875 26.74 27.075 ;
 RECT 26.516 26.875 26.572 27.075 ;
 RECT 25.676 26.875 25.732 27.075 ;
 RECT 25.508 26.875 25.564 27.075 ;
 RECT 26.012 26.875 26.068 27.075 ;
 RECT 25.844 26.875 25.9 27.075 ;
 RECT 25.34 26.875 25.396 27.075 ;
 END
 END vss.gds2219
 PIN vss.gds2220
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.314 26.9905 31.37 27.1905 ;
 END
 END vss.gds2220
 PIN vss.gds2221
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 29.642 30.95 29.842 ;
 END
 END vss.gds2221
 PIN vss.gds2222
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 29.682 31.922 29.882 ;
 END
 END vss.gds2222
 PIN vss.gds2223
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 26.2765 31.922 26.4765 ;
 END
 END vss.gds2223
 PIN vss.gds2224
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 26.2765 33.198 26.4765 ;
 END
 END vss.gds2224
 PIN vss.gds2225
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.314 29.231 30.37 29.431 ;
 END
 END vss.gds2225
 PIN vss.gds2226
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.49 29.023 34.546 29.223 ;
 END
 END vss.gds2226
 PIN vss.gds2227
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 26.52 33.866 26.72 ;
 END
 END vss.gds2227
 PIN vss.gds2228
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 30.397 33.198 30.597 ;
 END
 END vss.gds2228
 PIN vss.gds2229
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 28.4415 32.214 28.6415 ;
 END
 END vss.gds2229
 PIN vss.gds2230
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 28.224 34.046 28.424 ;
 END
 END vss.gds2230
 PIN vss.gds2231
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 30.0685 34.366 30.2685 ;
 END
 END vss.gds2231
 PIN vss.gds2232
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 30.197 32.47 30.397 ;
 END
 END vss.gds2232
 PIN vss.gds2233
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 28.2885 30.71 28.4885 ;
 END
 END vss.gds2233
 PIN vss.gds2234
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 26.4595 30.95 26.6595 ;
 END
 END vss.gds2234
 PIN vss.gds2235
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 28.5025 32.894 28.7025 ;
 END
 END vss.gds2235
 PIN vss.gds2236
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 28.277 33.542 28.477 ;
 END
 END vss.gds2236
 PIN vss.gds2237
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 29.137 33.198 29.337 ;
 END
 END vss.gds2237
 PIN vss.gds2238
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 28.5025 31.55 28.7025 ;
 END
 END vss.gds2238
 PIN vss.gds2239
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 28.3975 34.886 28.5975 ;
 END
 END vss.gds2239
 PIN vss.gds2240
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 30.296 28.469 30.352 28.669 ;
 RECT 32.228 26.122 32.284 26.322 ;
 RECT 32.06 26.122 32.116 26.322 ;
 RECT 30.716 26.103 30.772 26.303 ;
 RECT 30.548 26.103 30.604 26.303 ;
 RECT 31.052 26.103 31.108 26.303 ;
 RECT 31.22 26.103 31.276 26.303 ;
 RECT 30.884 26.103 30.94 26.303 ;
 RECT 31.892 26.103 31.948 26.303 ;
 RECT 31.556 26.122 31.612 26.322 ;
 RECT 31.724 26.122 31.78 26.322 ;
 RECT 33.152 26.122 33.208 26.322 ;
 RECT 32.648 26.122 32.704 26.322 ;
 RECT 32.48 26.122 32.536 26.322 ;
 RECT 32.816 26.122 32.872 26.322 ;
 RECT 33.656 26.122 33.712 26.322 ;
 RECT 33.824 26.122 33.88 26.322 ;
 RECT 33.488 26.122 33.544 26.322 ;
 RECT 33.32 26.122 33.376 26.322 ;
 RECT 34.748 26.122 34.804 26.322 ;
 RECT 34.328 26.103 34.384 26.285 ;
 RECT 34.076 26.103 34.132 26.285 ;
 RECT 32.312 25.842 32.368 26.042 ;
 RECT 30.296 25.842 30.352 26.042 ;
 RECT 30.632 25.842 30.688 26.042 ;
 RECT 30.968 25.842 31.024 26.042 ;
 RECT 31.304 25.842 31.36 26.042 ;
 RECT 31.976 25.842 32.032 26.042 ;
 RECT 32.648 25.842 32.704 26.042 ;
 RECT 32.984 25.842 33.04 26.042 ;
 RECT 33.32 25.842 33.376 26.042 ;
 RECT 34.244 25.879 34.3 26.061 ;
 RECT 33.992 25.879 34.048 26.061 ;
 RECT 34.58 25.842 34.636 26.042 ;
 RECT 34.832 25.842 34.888 26.042 ;
 RECT 32.648 28.804 32.704 29.004 ;
 RECT 32.9 28.807 32.956 29.007 ;
 RECT 33.572 29.84 33.628 29.993 ;
 RECT 31.052 29.82 31.108 29.993 ;
 RECT 31.22 29.793 31.276 29.993 ;
 RECT 32.816 29.837 32.872 30.002 ;
 RECT 32.648 29.837 32.704 30.002 ;
 RECT 31.892 29.837 31.948 30.002 ;
 RECT 31.724 29.837 31.78 30.002 ;
 RECT 32.648 30.064 32.704 30.264 ;
 RECT 32.9 30.067 32.956 30.267 ;
 RECT 35.168 26.654 35.224 26.854 ;
 RECT 31.388 30.413 31.444 30.613 ;
 RECT 31.22 30.413 31.276 30.613 ;
 RECT 30.464 27.673 30.52 27.873 ;
 RECT 32.06 29.363 32.116 29.563 ;
 RECT 32.48 29.363 32.536 29.563 ;
 RECT 31.388 29.153 31.444 29.353 ;
 RECT 31.22 29.153 31.276 29.353 ;
 RECT 30.716 29.287 30.772 29.487 ;
 RECT 33.404 29.4635 33.46 29.6635 ;
 RECT 33.908 29.2115 33.964 29.4115 ;
 END
 END vss.gds2240
 PIN vss.gds2241
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.698 25.982 39.738 26.182 ;
 END
 END vss.gds2241
 PIN vss.gds2242
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.026 25.982 39.066 26.182 ;
 END
 END vss.gds2242
 PIN vss.gds2243
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.354 25.982 38.394 26.182 ;
 END
 END vss.gds2243
 PIN vss.gds2244
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.682 25.982 37.722 26.182 ;
 END
 END vss.gds2244
 PIN vss.gds2245
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.01 25.982 37.05 26.182 ;
 END
 END vss.gds2245
 PIN vss.gds2246
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.338 25.982 36.378 26.182 ;
 END
 END vss.gds2246
 PIN vss.gds2247
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.666 25.982 35.706 26.182 ;
 END
 END vss.gds2247
 PIN vss.gds2248
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.102 25.775 40.148 25.975 ;
 END
 END vss.gds2248
 PIN vss.gds2249
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.43 25.775 39.476 25.975 ;
 END
 END vss.gds2249
 PIN vss.gds2250
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.826 25.775 39.866 25.975 ;
 END
 END vss.gds2250
 PIN vss.gds2251
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.758 25.775 38.804 25.975 ;
 END
 END vss.gds2251
 PIN vss.gds2252
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.154 25.775 39.194 25.975 ;
 END
 END vss.gds2252
 PIN vss.gds2253
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.086 25.775 38.132 25.975 ;
 END
 END vss.gds2253
 PIN vss.gds2254
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.482 25.775 38.522 25.975 ;
 END
 END vss.gds2254
 PIN vss.gds2255
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.414 25.775 37.46 25.975 ;
 END
 END vss.gds2255
 PIN vss.gds2256
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.81 25.775 37.85 25.975 ;
 END
 END vss.gds2256
 PIN vss.gds2257
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.742 25.775 36.788 25.975 ;
 END
 END vss.gds2257
 PIN vss.gds2258
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.138 25.775 37.178 25.975 ;
 END
 END vss.gds2258
 PIN vss.gds2259
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.07 25.775 36.116 25.975 ;
 END
 END vss.gds2259
 PIN vss.gds2260
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.466 25.775 36.506 25.975 ;
 END
 END vss.gds2260
 PIN vss.gds2261
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.398 25.775 35.444 25.975 ;
 END
 END vss.gds2261
 PIN vss.gds2262
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.794 25.775 35.834 25.975 ;
 END
 END vss.gds2262
 PIN vss.gds2263
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 28.2535 36.654 28.4535 ;
 END
 END vss.gds2263
 PIN vss.gds2264
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 28.2535 37.326 28.4535 ;
 END
 END vss.gds2264
 PIN vss.gds2265
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 28.2535 37.998 28.4535 ;
 END
 END vss.gds2265
 PIN vss.gds2266
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 28.2535 38.67 28.4535 ;
 END
 END vss.gds2266
 PIN vss.gds2267
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 28.2535 35.982 28.4535 ;
 END
 END vss.gds2267
 PIN vss.gds2268
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 28.2535 40.014 28.4535 ;
 END
 END vss.gds2268
 PIN vss.gds2269
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 27.837 35.31 28.037 ;
 END
 END vss.gds2269
 PIN vss.gds2270
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 28.2535 39.342 28.4535 ;
 END
 END vss.gds2270
 PIN vss.gds2271
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 39.956 28.563 40.012 28.763 ;
 RECT 39.788 28.573 39.844 28.773 ;
 RECT 39.284 28.563 39.34 28.763 ;
 RECT 39.116 28.573 39.172 28.773 ;
 RECT 38.612 28.563 38.668 28.763 ;
 RECT 38.444 28.573 38.5 28.773 ;
 RECT 37.94 28.563 37.996 28.763 ;
 RECT 37.772 28.573 37.828 28.773 ;
 RECT 37.268 28.563 37.324 28.763 ;
 RECT 37.1 28.573 37.156 28.773 ;
 RECT 36.596 28.563 36.652 28.763 ;
 RECT 36.428 28.573 36.484 28.773 ;
 RECT 35.252 28.563 35.308 28.763 ;
 RECT 35.924 28.563 35.98 28.763 ;
 RECT 35.756 28.573 35.812 28.773 ;
 RECT 39.62 25.801 39.676 26.001 ;
 RECT 39.452 25.801 39.508 26.001 ;
 RECT 39.788 25.816 39.844 26.016 ;
 RECT 39.956 25.816 40.012 26.016 ;
 RECT 38.948 25.801 39.004 26.001 ;
 RECT 38.78 25.801 38.836 26.001 ;
 RECT 39.116 25.816 39.172 26.016 ;
 RECT 39.284 25.816 39.34 26.016 ;
 RECT 38.276 25.801 38.332 26.001 ;
 RECT 38.108 25.801 38.164 26.001 ;
 RECT 38.444 25.816 38.5 26.016 ;
 RECT 38.612 25.816 38.668 26.016 ;
 RECT 37.604 25.801 37.66 26.001 ;
 RECT 37.436 25.801 37.492 26.001 ;
 RECT 37.772 25.816 37.828 26.016 ;
 RECT 37.94 25.816 37.996 26.016 ;
 RECT 36.932 25.801 36.988 26.001 ;
 RECT 36.764 25.801 36.82 26.001 ;
 RECT 37.1 25.816 37.156 26.016 ;
 RECT 37.268 25.816 37.324 26.016 ;
 RECT 36.26 25.801 36.316 26.001 ;
 RECT 36.092 25.801 36.148 26.001 ;
 RECT 36.428 25.816 36.484 26.016 ;
 RECT 36.596 25.816 36.652 26.016 ;
 RECT 35.252 25.816 35.308 26.016 ;
 RECT 35.756 25.816 35.812 26.016 ;
 RECT 35.924 25.816 35.98 26.016 ;
 RECT 40.124 25.801 40.18 26.001 ;
 RECT 35.588 25.801 35.644 26.001 ;
 RECT 35.42 25.801 35.476 26.001 ;
 RECT 40.124 26.875 40.18 27.075 ;
 RECT 39.62 26.875 39.676 27.075 ;
 RECT 39.452 26.875 39.508 27.075 ;
 RECT 39.956 26.875 40.012 27.075 ;
 RECT 39.788 26.875 39.844 27.075 ;
 RECT 38.948 26.875 39.004 27.075 ;
 RECT 38.78 26.875 38.836 27.075 ;
 RECT 39.284 26.875 39.34 27.075 ;
 RECT 39.116 26.875 39.172 27.075 ;
 RECT 38.276 26.875 38.332 27.075 ;
 RECT 38.108 26.875 38.164 27.075 ;
 RECT 38.612 26.875 38.668 27.075 ;
 RECT 38.444 26.875 38.5 27.075 ;
 RECT 37.604 26.875 37.66 27.075 ;
 RECT 37.436 26.875 37.492 27.075 ;
 RECT 37.94 26.875 37.996 27.075 ;
 RECT 37.772 26.875 37.828 27.075 ;
 RECT 36.932 26.875 36.988 27.075 ;
 RECT 36.764 26.875 36.82 27.075 ;
 RECT 37.268 26.875 37.324 27.075 ;
 RECT 37.1 26.875 37.156 27.075 ;
 RECT 36.26 26.875 36.316 27.075 ;
 RECT 36.092 26.875 36.148 27.075 ;
 RECT 36.596 26.875 36.652 27.075 ;
 RECT 36.428 26.875 36.484 27.075 ;
 RECT 35.588 26.875 35.644 27.075 ;
 RECT 35.252 26.875 35.308 27.075 ;
 RECT 35.42 26.875 35.476 27.075 ;
 RECT 35.924 26.875 35.98 27.075 ;
 RECT 35.756 26.875 35.812 27.075 ;
 END
 END vss.gds2271
 PIN vss.gds2272
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.822 25.982 44.862 26.182 ;
 END
 END vss.gds2272
 PIN vss.gds2273
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.15 25.982 44.19 26.182 ;
 END
 END vss.gds2273
 PIN vss.gds2274
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.478 25.982 43.518 26.182 ;
 END
 END vss.gds2274
 PIN vss.gds2275
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.806 25.982 42.846 26.182 ;
 END
 END vss.gds2275
 PIN vss.gds2276
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.134 25.982 42.174 26.182 ;
 END
 END vss.gds2276
 PIN vss.gds2277
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.462 25.982 41.502 26.182 ;
 END
 END vss.gds2277
 PIN vss.gds2278
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.37 25.982 40.41 26.182 ;
 END
 END vss.gds2278
 PIN vss.gds2279
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.226 25.775 45.272 25.975 ;
 END
 END vss.gds2279
 PIN vss.gds2280
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.554 25.775 44.6 25.975 ;
 END
 END vss.gds2280
 PIN vss.gds2281
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.95 25.775 44.99 25.975 ;
 END
 END vss.gds2281
 PIN vss.gds2282
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.882 25.775 43.928 25.975 ;
 END
 END vss.gds2282
 PIN vss.gds2283
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.278 25.775 44.318 25.975 ;
 END
 END vss.gds2283
 PIN vss.gds2284
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.21 25.775 43.256 25.975 ;
 END
 END vss.gds2284
 PIN vss.gds2285
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.606 25.775 43.646 25.975 ;
 END
 END vss.gds2285
 PIN vss.gds2286
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.538 25.775 42.584 25.975 ;
 END
 END vss.gds2286
 PIN vss.gds2287
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.934 25.775 42.974 25.975 ;
 END
 END vss.gds2287
 PIN vss.gds2288
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.866 25.775 41.912 25.975 ;
 END
 END vss.gds2288
 PIN vss.gds2289
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.262 25.775 42.302 25.975 ;
 END
 END vss.gds2289
 PIN vss.gds2290
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.194 25.775 41.24 25.975 ;
 END
 END vss.gds2290
 PIN vss.gds2291
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.59 25.775 41.63 25.975 ;
 END
 END vss.gds2291
 PIN vss.gds2292
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.498 25.775 40.538 25.975 ;
 END
 END vss.gds2292
 PIN vss.gds2293
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.774 26.9905 40.814 27.1905 ;
 END
 END vss.gds2293
 PIN vss.gds2294
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.918 26.9905 40.958 27.1905 ;
 END
 END vss.gds2294
 PIN vss.gds2295
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 28.2535 45.138 28.4535 ;
 END
 END vss.gds2295
 PIN vss.gds2296
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 28.2535 44.466 28.4535 ;
 END
 END vss.gds2296
 PIN vss.gds2297
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 28.2535 43.794 28.4535 ;
 END
 END vss.gds2297
 PIN vss.gds2298
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 28.2535 43.122 28.4535 ;
 END
 END vss.gds2298
 PIN vss.gds2299
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 28.2535 42.45 28.4535 ;
 END
 END vss.gds2299
 PIN vss.gds2300
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 28.2535 41.778 28.4535 ;
 END
 END vss.gds2300
 PIN vss.gds2301
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 28.2535 40.686 28.4535 ;
 END
 END vss.gds2301
 PIN vss.gds2302
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.046 26.9135 41.106 27.1135 ;
 END
 END vss.gds2302
 PIN vss.gds2303
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 45.08 28.563 45.136 28.763 ;
 RECT 44.912 28.573 44.968 28.773 ;
 RECT 44.408 28.563 44.464 28.763 ;
 RECT 44.24 28.573 44.296 28.773 ;
 RECT 43.736 28.563 43.792 28.763 ;
 RECT 43.568 28.573 43.624 28.773 ;
 RECT 43.064 28.563 43.12 28.763 ;
 RECT 42.896 28.573 42.952 28.773 ;
 RECT 42.392 28.563 42.448 28.763 ;
 RECT 42.224 28.573 42.28 28.773 ;
 RECT 41.048 28.563 41.104 28.763 ;
 RECT 41.72 28.563 41.776 28.763 ;
 RECT 41.552 28.573 41.608 28.773 ;
 RECT 40.628 28.563 40.684 28.763 ;
 RECT 40.46 28.573 40.516 28.773 ;
 RECT 44.744 25.801 44.8 26.001 ;
 RECT 44.576 25.801 44.632 26.001 ;
 RECT 44.912 25.816 44.968 26.016 ;
 RECT 45.08 25.816 45.136 26.016 ;
 RECT 44.072 25.801 44.128 26.001 ;
 RECT 43.904 25.801 43.96 26.001 ;
 RECT 44.24 25.816 44.296 26.016 ;
 RECT 44.408 25.816 44.464 26.016 ;
 RECT 43.4 25.801 43.456 26.001 ;
 RECT 43.232 25.801 43.288 26.001 ;
 RECT 43.568 25.816 43.624 26.016 ;
 RECT 43.736 25.816 43.792 26.016 ;
 RECT 42.728 25.801 42.784 26.001 ;
 RECT 42.56 25.801 42.616 26.001 ;
 RECT 42.896 25.816 42.952 26.016 ;
 RECT 43.064 25.816 43.12 26.016 ;
 RECT 42.056 25.801 42.112 26.001 ;
 RECT 41.888 25.801 41.944 26.001 ;
 RECT 42.224 25.816 42.28 26.016 ;
 RECT 42.392 25.816 42.448 26.016 ;
 RECT 41.048 25.816 41.104 26.016 ;
 RECT 41.552 25.816 41.608 26.016 ;
 RECT 41.72 25.816 41.776 26.016 ;
 RECT 40.46 25.816 40.516 26.016 ;
 RECT 40.628 25.816 40.684 26.016 ;
 RECT 41.384 25.801 41.44 26.001 ;
 RECT 41.216 25.801 41.272 26.001 ;
 RECT 40.292 25.801 40.348 26.001 ;
 RECT 40.964 29.3 41.02 29.5 ;
 RECT 44.744 26.875 44.8 27.075 ;
 RECT 44.576 26.875 44.632 27.075 ;
 RECT 45.08 26.875 45.136 27.075 ;
 RECT 44.912 26.875 44.968 27.075 ;
 RECT 44.072 26.875 44.128 27.075 ;
 RECT 43.904 26.875 43.96 27.075 ;
 RECT 44.408 26.875 44.464 27.075 ;
 RECT 44.24 26.875 44.296 27.075 ;
 RECT 43.4 26.875 43.456 27.075 ;
 RECT 43.232 26.875 43.288 27.075 ;
 RECT 43.736 26.875 43.792 27.075 ;
 RECT 43.568 26.875 43.624 27.075 ;
 RECT 42.728 26.875 42.784 27.075 ;
 RECT 42.56 26.875 42.616 27.075 ;
 RECT 43.064 26.875 43.12 27.075 ;
 RECT 42.896 26.875 42.952 27.075 ;
 RECT 42.056 26.875 42.112 27.075 ;
 RECT 41.888 26.875 41.944 27.075 ;
 RECT 42.392 26.875 42.448 27.075 ;
 RECT 42.224 26.875 42.28 27.075 ;
 RECT 41.384 26.875 41.44 27.075 ;
 RECT 41.048 26.875 41.104 27.075 ;
 RECT 41.216 26.875 41.272 27.075 ;
 RECT 41.72 26.875 41.776 27.075 ;
 RECT 41.552 26.875 41.608 27.075 ;
 RECT 40.628 26.875 40.684 27.075 ;
 RECT 40.46 26.875 40.516 27.075 ;
 RECT 40.292 26.875 40.348 27.075 ;
 RECT 40.796 28.7285 40.852 28.9285 ;
 END
 END vss.gds2303
 PIN vss.gds2304
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.366 26.9905 48.422 27.1905 ;
 END
 END vss.gds2304
 PIN vss.gds2305
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 29.642 48.002 29.842 ;
 END
 END vss.gds2305
 PIN vss.gds2306
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 29.682 48.974 29.882 ;
 END
 END vss.gds2306
 PIN vss.gds2307
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.166 25.982 46.206 26.182 ;
 END
 END vss.gds2307
 PIN vss.gds2308
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.494 25.982 45.534 26.182 ;
 END
 END vss.gds2308
 PIN vss.gds2309
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 26.2765 48.974 26.4765 ;
 END
 END vss.gds2309
 PIN vss.gds2310
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 26.2765 50.25 26.4765 ;
 END
 END vss.gds2310
 PIN vss.gds2311
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.898 25.775 45.944 25.975 ;
 END
 END vss.gds2311
 PIN vss.gds2312
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.294 25.775 46.334 25.975 ;
 END
 END vss.gds2312
 PIN vss.gds2313
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.622 25.775 45.662 25.975 ;
 END
 END vss.gds2313
 PIN vss.gds2314
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.366 29.231 47.422 29.431 ;
 END
 END vss.gds2314
 PIN vss.gds2315
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 27.837 46.482 28.037 ;
 END
 END vss.gds2315
 PIN vss.gds2316
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 28.2535 45.81 28.4535 ;
 END
 END vss.gds2316
 PIN vss.gds2317
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 26.102 47.162 26.302 ;
 END
 END vss.gds2317
 PIN vss.gds2318
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 30.197 49.522 30.397 ;
 END
 END vss.gds2318
 PIN vss.gds2319
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 28.3975 46.922 28.5975 ;
 END
 END vss.gds2319
 PIN vss.gds2320
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 26.4595 48.002 26.6595 ;
 END
 END vss.gds2320
 PIN vss.gds2321
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 27.6625 46.694 27.8625 ;
 END
 END vss.gds2321
 PIN vss.gds2322
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 28.2885 47.762 28.4885 ;
 END
 END vss.gds2322
 PIN vss.gds2323
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 28.4415 49.266 28.6415 ;
 END
 END vss.gds2323
 PIN vss.gds2324
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 30.397 50.25 30.597 ;
 END
 END vss.gds2324
 PIN vss.gds2325
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 29.137 50.25 29.337 ;
 END
 END vss.gds2325
 PIN vss.gds2326
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 28.5025 48.602 28.7025 ;
 END
 END vss.gds2326
 PIN vss.gds2327
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 28.5025 49.946 28.7025 ;
 END
 END vss.gds2327
 PIN vss.gds2328
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 47.348 28.469 47.404 28.669 ;
 RECT 46.424 28.563 46.48 28.763 ;
 RECT 46.256 28.573 46.312 28.773 ;
 RECT 45.752 28.563 45.808 28.763 ;
 RECT 45.584 28.573 45.64 28.773 ;
 RECT 46.928 26.122 46.984 26.322 ;
 RECT 49.28 26.122 49.336 26.322 ;
 RECT 49.112 26.122 49.168 26.322 ;
 RECT 47.768 26.103 47.824 26.303 ;
 RECT 47.096 26.103 47.152 26.303 ;
 RECT 47.264 26.103 47.32 26.303 ;
 RECT 47.6 26.103 47.656 26.303 ;
 RECT 48.104 26.103 48.16 26.303 ;
 RECT 48.272 26.103 48.328 26.303 ;
 RECT 47.936 26.103 47.992 26.303 ;
 RECT 48.944 26.103 49 26.303 ;
 RECT 48.608 26.122 48.664 26.322 ;
 RECT 48.776 26.122 48.832 26.322 ;
 RECT 50.204 26.122 50.26 26.322 ;
 RECT 49.7 26.122 49.756 26.322 ;
 RECT 49.532 26.122 49.588 26.322 ;
 RECT 49.868 26.122 49.924 26.322 ;
 RECT 49.364 25.842 49.42 26.042 ;
 RECT 47.348 25.842 47.404 26.042 ;
 RECT 47.684 25.842 47.74 26.042 ;
 RECT 47.012 25.842 47.068 26.042 ;
 RECT 48.02 25.842 48.076 26.042 ;
 RECT 48.356 25.842 48.412 26.042 ;
 RECT 49.028 25.842 49.084 26.042 ;
 RECT 49.7 25.842 49.756 26.042 ;
 RECT 50.036 25.842 50.092 26.042 ;
 RECT 46.088 25.801 46.144 26.001 ;
 RECT 45.92 25.801 45.976 26.001 ;
 RECT 46.256 25.816 46.312 26.016 ;
 RECT 46.424 25.816 46.48 26.016 ;
 RECT 45.416 25.801 45.472 26.001 ;
 RECT 45.248 25.801 45.304 26.001 ;
 RECT 45.584 25.816 45.64 26.016 ;
 RECT 45.752 25.816 45.808 26.016 ;
 RECT 49.7 28.804 49.756 29.004 ;
 RECT 49.952 28.807 50.008 29.007 ;
 RECT 48.104 29.82 48.16 29.993 ;
 RECT 48.272 29.793 48.328 29.993 ;
 RECT 49.868 29.837 49.924 30.002 ;
 RECT 49.7 29.837 49.756 30.002 ;
 RECT 48.944 29.837 49 30.002 ;
 RECT 48.776 29.837 48.832 30.002 ;
 RECT 49.7 30.064 49.756 30.264 ;
 RECT 49.952 30.067 50.008 30.267 ;
 RECT 47.264 27.459 47.32 27.659 ;
 RECT 47.516 27.673 47.572 27.873 ;
 RECT 48.44 30.413 48.496 30.613 ;
 RECT 48.272 30.413 48.328 30.613 ;
 RECT 49.112 29.363 49.168 29.563 ;
 RECT 49.532 29.363 49.588 29.563 ;
 RECT 48.44 29.153 48.496 29.353 ;
 RECT 48.272 29.153 48.328 29.353 ;
 RECT 47.768 29.287 47.824 29.487 ;
 RECT 46.088 26.875 46.144 27.075 ;
 RECT 45.92 26.875 45.976 27.075 ;
 RECT 46.424 26.875 46.48 27.075 ;
 RECT 46.256 26.875 46.312 27.075 ;
 RECT 45.416 26.875 45.472 27.075 ;
 RECT 45.248 26.875 45.304 27.075 ;
 RECT 45.752 26.875 45.808 27.075 ;
 RECT 45.584 26.875 45.64 27.075 ;
 END
 END vss.gds2328
 PIN vss.gds2329
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.734 25.982 54.774 26.182 ;
 END
 END vss.gds2329
 PIN vss.gds2330
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.062 25.982 54.102 26.182 ;
 END
 END vss.gds2330
 PIN vss.gds2331
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.39 25.982 53.43 26.182 ;
 END
 END vss.gds2331
 PIN vss.gds2332
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.718 25.982 52.758 26.182 ;
 END
 END vss.gds2332
 PIN vss.gds2333
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.138 25.775 55.184 25.975 ;
 END
 END vss.gds2333
 PIN vss.gds2334
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.466 25.775 54.512 25.975 ;
 END
 END vss.gds2334
 PIN vss.gds2335
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.862 25.775 54.902 25.975 ;
 END
 END vss.gds2335
 PIN vss.gds2336
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.794 25.775 53.84 25.975 ;
 END
 END vss.gds2336
 PIN vss.gds2337
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.19 25.775 54.23 25.975 ;
 END
 END vss.gds2337
 PIN vss.gds2338
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.122 25.775 53.168 25.975 ;
 END
 END vss.gds2338
 PIN vss.gds2339
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.518 25.775 53.558 25.975 ;
 END
 END vss.gds2339
 PIN vss.gds2340
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.45 25.775 52.496 25.975 ;
 END
 END vss.gds2340
 PIN vss.gds2341
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.846 25.775 52.886 25.975 ;
 END
 END vss.gds2341
 PIN vss.gds2342
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.542 29.023 51.598 29.223 ;
 END
 END vss.gds2342
 PIN vss.gds2343
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 26.52 50.918 26.72 ;
 END
 END vss.gds2343
 PIN vss.gds2344
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 28.2535 55.05 28.4535 ;
 END
 END vss.gds2344
 PIN vss.gds2345
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 28.2535 54.378 28.4535 ;
 END
 END vss.gds2345
 PIN vss.gds2346
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 28.2535 53.706 28.4535 ;
 END
 END vss.gds2346
 PIN vss.gds2347
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 30.0685 51.418 30.2685 ;
 END
 END vss.gds2347
 PIN vss.gds2348
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 28.224 51.098 28.424 ;
 END
 END vss.gds2348
 PIN vss.gds2349
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 28.2535 53.034 28.4535 ;
 END
 END vss.gds2349
 PIN vss.gds2350
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 28.3975 51.938 28.5975 ;
 END
 END vss.gds2350
 PIN vss.gds2351
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 28.277 50.594 28.477 ;
 END
 END vss.gds2351
 PIN vss.gds2352
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 27.837 52.362 28.037 ;
 END
 END vss.gds2352
 PIN vss.gds2353
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 54.992 28.563 55.048 28.763 ;
 RECT 54.824 28.573 54.88 28.773 ;
 RECT 54.32 28.563 54.376 28.763 ;
 RECT 54.152 28.573 54.208 28.773 ;
 RECT 53.648 28.563 53.704 28.763 ;
 RECT 53.48 28.573 53.536 28.773 ;
 RECT 52.304 28.563 52.36 28.763 ;
 RECT 52.976 28.563 53.032 28.763 ;
 RECT 52.808 28.573 52.864 28.773 ;
 RECT 50.708 26.122 50.764 26.322 ;
 RECT 50.876 26.122 50.932 26.322 ;
 RECT 50.54 26.122 50.596 26.322 ;
 RECT 50.372 26.122 50.428 26.322 ;
 RECT 51.8 26.122 51.856 26.322 ;
 RECT 51.38 26.103 51.436 26.285 ;
 RECT 51.128 26.103 51.184 26.285 ;
 RECT 55.16 25.801 55.216 26.001 ;
 RECT 54.656 25.801 54.712 26.001 ;
 RECT 54.488 25.801 54.544 26.001 ;
 RECT 54.824 25.816 54.88 26.016 ;
 RECT 54.992 25.816 55.048 26.016 ;
 RECT 53.984 25.801 54.04 26.001 ;
 RECT 53.816 25.801 53.872 26.001 ;
 RECT 54.152 25.816 54.208 26.016 ;
 RECT 54.32 25.816 54.376 26.016 ;
 RECT 50.372 25.842 50.428 26.042 ;
 RECT 51.296 25.879 51.352 26.061 ;
 RECT 51.044 25.879 51.1 26.061 ;
 RECT 51.632 25.842 51.688 26.042 ;
 RECT 51.884 25.842 51.94 26.042 ;
 RECT 53.312 25.801 53.368 26.001 ;
 RECT 53.144 25.801 53.2 26.001 ;
 RECT 53.48 25.816 53.536 26.016 ;
 RECT 53.648 25.816 53.704 26.016 ;
 RECT 52.304 25.816 52.36 26.016 ;
 RECT 52.808 25.816 52.864 26.016 ;
 RECT 52.976 25.816 53.032 26.016 ;
 RECT 50.624 29.84 50.68 29.993 ;
 RECT 52.64 25.801 52.696 26.001 ;
 RECT 52.472 25.801 52.528 26.001 ;
 RECT 52.22 26.654 52.276 26.854 ;
 RECT 50.96 29.2115 51.016 29.4115 ;
 RECT 50.456 29.4635 50.512 29.6635 ;
 RECT 55.16 26.875 55.216 27.075 ;
 RECT 54.656 26.875 54.712 27.075 ;
 RECT 54.488 26.875 54.544 27.075 ;
 RECT 54.992 26.875 55.048 27.075 ;
 RECT 54.824 26.875 54.88 27.075 ;
 RECT 53.984 26.875 54.04 27.075 ;
 RECT 53.816 26.875 53.872 27.075 ;
 RECT 54.32 26.875 54.376 27.075 ;
 RECT 54.152 26.875 54.208 27.075 ;
 RECT 53.312 26.875 53.368 27.075 ;
 RECT 53.144 26.875 53.2 27.075 ;
 RECT 53.648 26.875 53.704 27.075 ;
 RECT 53.48 26.875 53.536 27.075 ;
 RECT 52.64 26.875 52.696 27.075 ;
 RECT 52.304 26.875 52.36 27.075 ;
 RECT 52.472 26.875 52.528 27.075 ;
 RECT 52.976 26.875 53.032 27.075 ;
 RECT 52.808 26.875 52.864 27.075 ;
 END
 END vss.gds2353
 PIN vss.gds2354
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.858 25.982 59.898 26.182 ;
 END
 END vss.gds2354
 PIN vss.gds2355
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.186 25.982 59.226 26.182 ;
 END
 END vss.gds2355
 PIN vss.gds2356
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.514 25.982 58.554 26.182 ;
 END
 END vss.gds2356
 PIN vss.gds2357
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.422 25.982 57.462 26.182 ;
 END
 END vss.gds2357
 PIN vss.gds2358
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.75 25.982 56.79 26.182 ;
 END
 END vss.gds2358
 PIN vss.gds2359
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.078 25.982 56.118 26.182 ;
 END
 END vss.gds2359
 PIN vss.gds2360
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.406 25.982 55.446 26.182 ;
 END
 END vss.gds2360
 PIN vss.gds2361
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.59 25.775 59.636 25.975 ;
 END
 END vss.gds2361
 PIN vss.gds2362
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.986 25.775 60.026 25.975 ;
 END
 END vss.gds2362
 PIN vss.gds2363
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.918 25.775 58.964 25.975 ;
 END
 END vss.gds2363
 PIN vss.gds2364
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.314 25.775 59.354 25.975 ;
 END
 END vss.gds2364
 PIN vss.gds2365
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.246 25.775 58.292 25.975 ;
 END
 END vss.gds2365
 PIN vss.gds2366
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.642 25.775 58.682 25.975 ;
 END
 END vss.gds2366
 PIN vss.gds2367
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.154 25.775 57.2 25.975 ;
 END
 END vss.gds2367
 PIN vss.gds2368
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.55 25.775 57.59 25.975 ;
 END
 END vss.gds2368
 PIN vss.gds2369
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.482 25.775 56.528 25.975 ;
 END
 END vss.gds2369
 PIN vss.gds2370
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.878 25.775 56.918 25.975 ;
 END
 END vss.gds2370
 PIN vss.gds2371
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.81 25.775 55.856 25.975 ;
 END
 END vss.gds2371
 PIN vss.gds2372
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.206 25.775 56.246 25.975 ;
 END
 END vss.gds2372
 PIN vss.gds2373
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.534 25.775 55.574 25.975 ;
 END
 END vss.gds2373
 PIN vss.gds2374
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.826 26.9905 57.866 27.1905 ;
 END
 END vss.gds2374
 PIN vss.gds2375
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.97 26.9905 58.01 27.1905 ;
 END
 END vss.gds2375
 PIN vss.gds2376
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.098 26.9135 58.158 27.1135 ;
 END
 END vss.gds2376
 PIN vss.gds2377
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 28.2535 60.174 28.4535 ;
 END
 END vss.gds2377
 PIN vss.gds2378
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 28.2535 59.502 28.4535 ;
 END
 END vss.gds2378
 PIN vss.gds2379
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 28.2535 58.83 28.4535 ;
 END
 END vss.gds2379
 PIN vss.gds2380
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 28.2535 55.722 28.4535 ;
 END
 END vss.gds2380
 PIN vss.gds2381
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 28.2535 56.394 28.4535 ;
 END
 END vss.gds2381
 PIN vss.gds2382
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 28.2535 57.738 28.4535 ;
 END
 END vss.gds2382
 PIN vss.gds2383
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 28.2535 57.066 28.4535 ;
 END
 END vss.gds2383
 PIN vss.gds2384
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 60.116 28.563 60.172 28.763 ;
 RECT 59.948 28.573 60.004 28.773 ;
 RECT 59.444 28.563 59.5 28.763 ;
 RECT 59.276 28.573 59.332 28.773 ;
 RECT 58.1 28.563 58.156 28.763 ;
 RECT 58.772 28.563 58.828 28.763 ;
 RECT 58.604 28.573 58.66 28.773 ;
 RECT 57.68 28.563 57.736 28.763 ;
 RECT 57.512 28.573 57.568 28.773 ;
 RECT 57.008 28.563 57.064 28.763 ;
 RECT 56.84 28.573 56.896 28.773 ;
 RECT 56.336 28.563 56.392 28.763 ;
 RECT 56.168 28.573 56.224 28.773 ;
 RECT 55.664 28.563 55.72 28.763 ;
 RECT 55.496 28.573 55.552 28.773 ;
 RECT 59.78 25.801 59.836 26.001 ;
 RECT 59.612 25.801 59.668 26.001 ;
 RECT 59.948 25.816 60.004 26.016 ;
 RECT 60.116 25.816 60.172 26.016 ;
 RECT 59.108 25.801 59.164 26.001 ;
 RECT 58.94 25.801 58.996 26.001 ;
 RECT 59.276 25.816 59.332 26.016 ;
 RECT 59.444 25.816 59.5 26.016 ;
 RECT 58.1 25.816 58.156 26.016 ;
 RECT 58.604 25.816 58.66 26.016 ;
 RECT 58.772 25.816 58.828 26.016 ;
 RECT 57.512 25.816 57.568 26.016 ;
 RECT 57.68 25.816 57.736 26.016 ;
 RECT 56.672 25.801 56.728 26.001 ;
 RECT 56.504 25.801 56.56 26.001 ;
 RECT 56.84 25.816 56.896 26.016 ;
 RECT 57.008 25.816 57.064 26.016 ;
 RECT 56 25.801 56.056 26.001 ;
 RECT 55.832 25.801 55.888 26.001 ;
 RECT 56.168 25.816 56.224 26.016 ;
 RECT 56.336 25.816 56.392 26.016 ;
 RECT 55.328 25.801 55.384 26.001 ;
 RECT 55.496 25.816 55.552 26.016 ;
 RECT 55.664 25.816 55.72 26.016 ;
 RECT 59.78 26.875 59.836 27.075 ;
 RECT 59.612 26.875 59.668 27.075 ;
 RECT 60.116 26.875 60.172 27.075 ;
 RECT 59.948 26.875 60.004 27.075 ;
 RECT 59.108 26.875 59.164 27.075 ;
 RECT 58.94 26.875 58.996 27.075 ;
 RECT 59.444 26.875 59.5 27.075 ;
 RECT 59.276 26.875 59.332 27.075 ;
 RECT 58.436 26.875 58.492 27.075 ;
 RECT 58.1 26.875 58.156 27.075 ;
 RECT 58.268 26.875 58.324 27.075 ;
 RECT 58.772 26.875 58.828 27.075 ;
 RECT 58.604 26.875 58.66 27.075 ;
 RECT 58.436 25.801 58.492 26.001 ;
 RECT 58.268 25.801 58.324 26.001 ;
 RECT 57.344 25.801 57.4 26.001 ;
 RECT 57.176 25.801 57.232 26.001 ;
 RECT 58.016 29.3 58.072 29.5 ;
 RECT 57.344 26.875 57.4 27.075 ;
 RECT 57.176 26.875 57.232 27.075 ;
 RECT 57.68 26.875 57.736 27.075 ;
 RECT 57.512 26.875 57.568 27.075 ;
 RECT 56.672 26.875 56.728 27.075 ;
 RECT 56.504 26.875 56.56 27.075 ;
 RECT 57.008 26.875 57.064 27.075 ;
 RECT 56.84 26.875 56.896 27.075 ;
 RECT 56 26.875 56.056 27.075 ;
 RECT 55.832 26.875 55.888 27.075 ;
 RECT 56.336 26.875 56.392 27.075 ;
 RECT 56.168 26.875 56.224 27.075 ;
 RECT 55.328 26.875 55.384 27.075 ;
 RECT 55.664 26.875 55.72 27.075 ;
 RECT 55.496 26.875 55.552 27.075 ;
 RECT 57.848 28.7285 57.904 28.9285 ;
 END
 END vss.gds2384
 PIN vss.gds2385
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 29.642 65.054 29.842 ;
 END
 END vss.gds2385
 PIN vss.gds2386
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.218 25.982 63.258 26.182 ;
 END
 END vss.gds2386
 PIN vss.gds2387
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.546 25.982 62.586 26.182 ;
 END
 END vss.gds2387
 PIN vss.gds2388
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.874 25.982 61.914 26.182 ;
 END
 END vss.gds2388
 PIN vss.gds2389
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.202 25.982 61.242 26.182 ;
 END
 END vss.gds2389
 PIN vss.gds2390
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.53 25.982 60.57 26.182 ;
 END
 END vss.gds2390
 PIN vss.gds2391
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.95 25.775 62.996 25.975 ;
 END
 END vss.gds2391
 PIN vss.gds2392
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.346 25.775 63.386 25.975 ;
 END
 END vss.gds2392
 PIN vss.gds2393
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.278 25.775 62.324 25.975 ;
 END
 END vss.gds2393
 PIN vss.gds2394
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.674 25.775 62.714 25.975 ;
 END
 END vss.gds2394
 PIN vss.gds2395
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.606 25.775 61.652 25.975 ;
 END
 END vss.gds2395
 PIN vss.gds2396
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.002 25.775 62.042 25.975 ;
 END
 END vss.gds2396
 PIN vss.gds2397
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.934 25.775 60.98 25.975 ;
 END
 END vss.gds2397
 PIN vss.gds2398
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.33 25.775 61.37 25.975 ;
 END
 END vss.gds2398
 PIN vss.gds2399
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.262 25.775 60.308 25.975 ;
 END
 END vss.gds2399
 PIN vss.gds2400
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.658 25.775 60.698 25.975 ;
 END
 END vss.gds2400
 PIN vss.gds2401
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 26.102 64.214 26.302 ;
 END
 END vss.gds2401
 PIN vss.gds2402
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.418 29.231 64.474 29.431 ;
 END
 END vss.gds2402
 PIN vss.gds2403
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 27.837 63.534 28.037 ;
 END
 END vss.gds2403
 PIN vss.gds2404
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 28.2535 62.862 28.4535 ;
 END
 END vss.gds2404
 PIN vss.gds2405
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 28.2535 62.19 28.4535 ;
 END
 END vss.gds2405
 PIN vss.gds2406
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 28.2535 61.518 28.4535 ;
 END
 END vss.gds2406
 PIN vss.gds2407
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 28.2535 60.846 28.4535 ;
 END
 END vss.gds2407
 PIN vss.gds2408
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 28.3975 63.974 28.5975 ;
 END
 END vss.gds2408
 PIN vss.gds2409
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 27.6625 63.746 27.8625 ;
 END
 END vss.gds2409
 PIN vss.gds2410
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 26.4595 65.054 26.6595 ;
 END
 END vss.gds2410
 PIN vss.gds2411
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 28.2885 64.814 28.4885 ;
 END
 END vss.gds2411
 PIN vss.gds2412
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 64.4 28.469 64.456 28.669 ;
 RECT 63.476 28.563 63.532 28.763 ;
 RECT 63.308 28.573 63.364 28.773 ;
 RECT 62.804 28.563 62.86 28.763 ;
 RECT 62.636 28.573 62.692 28.773 ;
 RECT 62.132 28.563 62.188 28.763 ;
 RECT 61.964 28.573 62.02 28.773 ;
 RECT 61.46 28.563 61.516 28.763 ;
 RECT 61.292 28.573 61.348 28.773 ;
 RECT 60.788 28.563 60.844 28.763 ;
 RECT 60.62 28.573 60.676 28.773 ;
 RECT 63.98 26.122 64.036 26.322 ;
 RECT 64.82 26.103 64.876 26.303 ;
 RECT 64.148 26.103 64.204 26.303 ;
 RECT 64.316 26.103 64.372 26.303 ;
 RECT 64.652 26.103 64.708 26.303 ;
 RECT 65.156 26.103 65.212 26.303 ;
 RECT 64.988 26.103 65.044 26.303 ;
 RECT 64.4 25.842 64.456 26.042 ;
 RECT 64.736 25.842 64.792 26.042 ;
 RECT 64.064 25.842 64.12 26.042 ;
 RECT 65.072 25.842 65.128 26.042 ;
 RECT 63.14 25.801 63.196 26.001 ;
 RECT 62.972 25.801 63.028 26.001 ;
 RECT 63.308 25.816 63.364 26.016 ;
 RECT 63.476 25.816 63.532 26.016 ;
 RECT 62.468 25.801 62.524 26.001 ;
 RECT 62.3 25.801 62.356 26.001 ;
 RECT 62.636 25.816 62.692 26.016 ;
 RECT 62.804 25.816 62.86 26.016 ;
 RECT 61.796 25.801 61.852 26.001 ;
 RECT 61.628 25.801 61.684 26.001 ;
 RECT 61.964 25.816 62.02 26.016 ;
 RECT 62.132 25.816 62.188 26.016 ;
 RECT 61.124 25.801 61.18 26.001 ;
 RECT 60.956 25.801 61.012 26.001 ;
 RECT 61.292 25.816 61.348 26.016 ;
 RECT 61.46 25.816 61.516 26.016 ;
 RECT 60.62 25.816 60.676 26.016 ;
 RECT 60.788 25.816 60.844 26.016 ;
 RECT 60.452 25.801 60.508 26.001 ;
 RECT 60.284 25.801 60.34 26.001 ;
 RECT 63.14 26.875 63.196 27.075 ;
 RECT 62.972 26.875 63.028 27.075 ;
 RECT 63.476 26.875 63.532 27.075 ;
 RECT 63.308 26.875 63.364 27.075 ;
 RECT 62.468 26.875 62.524 27.075 ;
 RECT 62.3 26.875 62.356 27.075 ;
 RECT 62.804 26.875 62.86 27.075 ;
 RECT 62.636 26.875 62.692 27.075 ;
 RECT 61.796 26.875 61.852 27.075 ;
 RECT 61.628 26.875 61.684 27.075 ;
 RECT 62.132 26.875 62.188 27.075 ;
 RECT 61.964 26.875 62.02 27.075 ;
 RECT 61.124 26.875 61.18 27.075 ;
 RECT 60.956 26.875 61.012 27.075 ;
 RECT 61.46 26.875 61.516 27.075 ;
 RECT 61.292 26.875 61.348 27.075 ;
 RECT 60.452 26.875 60.508 27.075 ;
 RECT 60.788 26.875 60.844 27.075 ;
 RECT 60.62 26.875 60.676 27.075 ;
 RECT 60.284 26.875 60.34 27.075 ;
 RECT 65.156 29.82 65.212 29.993 ;
 RECT 64.82 29.287 64.876 29.487 ;
 RECT 64.316 27.459 64.372 27.659 ;
 RECT 64.568 27.673 64.624 27.873 ;
 END
 END vss.gds2412
 PIN vss.gds2413
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.418 26.9905 65.474 27.1905 ;
 END
 END vss.gds2413
 PIN vss.gds2414
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 29.682 66.026 29.882 ;
 END
 END vss.gds2414
 PIN vss.gds2415
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.77 25.982 69.81 26.182 ;
 END
 END vss.gds2415
 PIN vss.gds2416
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 26.2765 66.026 26.4765 ;
 END
 END vss.gds2416
 PIN vss.gds2417
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 26.2765 67.302 26.4765 ;
 END
 END vss.gds2417
 PIN vss.gds2418
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.174 25.775 70.22 25.975 ;
 END
 END vss.gds2418
 PIN vss.gds2419
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.502 25.775 69.548 25.975 ;
 END
 END vss.gds2419
 PIN vss.gds2420
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.898 25.775 69.938 25.975 ;
 END
 END vss.gds2420
 PIN vss.gds2421
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 30.197 66.574 30.397 ;
 END
 END vss.gds2421
 PIN vss.gds2422
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.594 29.023 68.65 29.223 ;
 END
 END vss.gds2422
 PIN vss.gds2423
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 28.224 68.15 28.424 ;
 END
 END vss.gds2423
 PIN vss.gds2424
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 26.52 67.97 26.72 ;
 END
 END vss.gds2424
 PIN vss.gds2425
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 28.4415 66.318 28.6415 ;
 END
 END vss.gds2425
 PIN vss.gds2426
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 30.0685 68.47 30.2685 ;
 END
 END vss.gds2426
 PIN vss.gds2427
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 30.397 67.302 30.597 ;
 END
 END vss.gds2427
 PIN vss.gds2428
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 29.137 67.302 29.337 ;
 END
 END vss.gds2428
 PIN vss.gds2429
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 28.2535 70.086 28.4535 ;
 END
 END vss.gds2429
 PIN vss.gds2430
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 28.5025 66.998 28.7025 ;
 END
 END vss.gds2430
 PIN vss.gds2431
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 28.5025 65.654 28.7025 ;
 END
 END vss.gds2431
 PIN vss.gds2432
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 28.277 67.646 28.477 ;
 END
 END vss.gds2432
 PIN vss.gds2433
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 28.3975 68.99 28.5975 ;
 END
 END vss.gds2433
 PIN vss.gds2434
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 27.837 69.414 28.037 ;
 END
 END vss.gds2434
 PIN vss.gds2435
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 69.356 28.563 69.412 28.763 ;
 RECT 70.028 28.563 70.084 28.763 ;
 RECT 69.86 28.573 69.916 28.773 ;
 RECT 66.332 26.122 66.388 26.322 ;
 RECT 66.164 26.122 66.22 26.322 ;
 RECT 65.324 26.103 65.38 26.303 ;
 RECT 65.996 26.103 66.052 26.303 ;
 RECT 65.66 26.122 65.716 26.322 ;
 RECT 65.828 26.122 65.884 26.322 ;
 RECT 67.256 26.122 67.312 26.322 ;
 RECT 66.752 26.122 66.808 26.322 ;
 RECT 66.584 26.122 66.64 26.322 ;
 RECT 66.92 26.122 66.976 26.322 ;
 RECT 67.76 26.122 67.816 26.322 ;
 RECT 67.928 26.122 67.984 26.322 ;
 RECT 67.592 26.122 67.648 26.322 ;
 RECT 67.424 26.122 67.48 26.322 ;
 RECT 68.852 26.122 68.908 26.322 ;
 RECT 68.432 26.103 68.488 26.285 ;
 RECT 68.18 26.103 68.236 26.285 ;
 RECT 66.416 25.842 66.472 26.042 ;
 RECT 65.408 25.842 65.464 26.042 ;
 RECT 66.08 25.842 66.136 26.042 ;
 RECT 66.752 25.842 66.808 26.042 ;
 RECT 67.088 25.842 67.144 26.042 ;
 RECT 67.424 25.842 67.48 26.042 ;
 RECT 68.348 25.879 68.404 26.061 ;
 RECT 68.096 25.879 68.152 26.061 ;
 RECT 68.684 25.842 68.74 26.042 ;
 RECT 68.936 25.842 68.992 26.042 ;
 RECT 70.196 25.801 70.252 26.001 ;
 RECT 69.356 25.816 69.412 26.016 ;
 RECT 69.86 25.816 69.916 26.016 ;
 RECT 70.028 25.816 70.084 26.016 ;
 RECT 70.196 26.875 70.252 27.075 ;
 RECT 69.692 26.875 69.748 27.075 ;
 RECT 69.356 26.875 69.412 27.075 ;
 RECT 69.524 26.875 69.58 27.075 ;
 RECT 70.028 26.875 70.084 27.075 ;
 RECT 69.86 26.875 69.916 27.075 ;
 RECT 66.752 28.804 66.808 29.004 ;
 RECT 67.004 28.807 67.06 29.007 ;
 RECT 67.676 29.84 67.732 29.993 ;
 RECT 65.324 29.793 65.38 29.993 ;
 RECT 66.92 29.837 66.976 30.002 ;
 RECT 66.752 29.837 66.808 30.002 ;
 RECT 65.996 29.837 66.052 30.002 ;
 RECT 65.828 29.837 65.884 30.002 ;
 RECT 65.492 29.153 65.548 29.353 ;
 RECT 65.324 29.153 65.38 29.353 ;
 RECT 69.692 25.801 69.748 26.001 ;
 RECT 69.524 25.801 69.58 26.001 ;
 RECT 66.752 30.064 66.808 30.264 ;
 RECT 67.004 30.067 67.06 30.267 ;
 RECT 69.272 26.654 69.328 26.854 ;
 RECT 65.492 30.413 65.548 30.613 ;
 RECT 65.324 30.413 65.38 30.613 ;
 RECT 66.164 29.363 66.22 29.563 ;
 RECT 66.584 29.363 66.64 29.563 ;
 RECT 67.508 29.4635 67.564 29.6635 ;
 RECT 68.012 29.2115 68.068 29.4115 ;
 END
 END vss.gds2435
 PIN vss.gds2436
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.474 25.982 74.514 26.182 ;
 END
 END vss.gds2436
 PIN vss.gds2437
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.802 25.982 73.842 26.182 ;
 END
 END vss.gds2437
 PIN vss.gds2438
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.13 25.982 73.17 26.182 ;
 END
 END vss.gds2438
 PIN vss.gds2439
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.458 25.982 72.498 26.182 ;
 END
 END vss.gds2439
 PIN vss.gds2440
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.786 25.982 71.826 26.182 ;
 END
 END vss.gds2440
 PIN vss.gds2441
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.114 25.982 71.154 26.182 ;
 END
 END vss.gds2441
 PIN vss.gds2442
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.442 25.982 70.482 26.182 ;
 END
 END vss.gds2442
 PIN vss.gds2443
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.206 25.775 74.252 25.975 ;
 END
 END vss.gds2443
 PIN vss.gds2444
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.602 25.775 74.642 25.975 ;
 END
 END vss.gds2444
 PIN vss.gds2445
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.534 25.775 73.58 25.975 ;
 END
 END vss.gds2445
 PIN vss.gds2446
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.93 25.775 73.97 25.975 ;
 END
 END vss.gds2446
 PIN vss.gds2447
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.862 25.775 72.908 25.975 ;
 END
 END vss.gds2447
 PIN vss.gds2448
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.258 25.775 73.298 25.975 ;
 END
 END vss.gds2448
 PIN vss.gds2449
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.19 25.775 72.236 25.975 ;
 END
 END vss.gds2449
 PIN vss.gds2450
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.586 25.775 72.626 25.975 ;
 END
 END vss.gds2450
 PIN vss.gds2451
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.518 25.775 71.564 25.975 ;
 END
 END vss.gds2451
 PIN vss.gds2452
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.914 25.775 71.954 25.975 ;
 END
 END vss.gds2452
 PIN vss.gds2453
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.846 25.775 70.892 25.975 ;
 END
 END vss.gds2453
 PIN vss.gds2454
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.242 25.775 71.282 25.975 ;
 END
 END vss.gds2454
 PIN vss.gds2455
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.57 25.775 70.61 25.975 ;
 END
 END vss.gds2455
 PIN vss.gds2456
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 28.2535 71.43 28.4535 ;
 END
 END vss.gds2456
 PIN vss.gds2457
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 28.2535 72.102 28.4535 ;
 END
 END vss.gds2457
 PIN vss.gds2458
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 28.2535 72.774 28.4535 ;
 END
 END vss.gds2458
 PIN vss.gds2459
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 28.2535 70.758 28.4535 ;
 END
 END vss.gds2459
 PIN vss.gds2460
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 28.2535 73.446 28.4535 ;
 END
 END vss.gds2460
 PIN vss.gds2461
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 28.2535 74.118 28.4535 ;
 END
 END vss.gds2461
 PIN vss.gds2462
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 28.2535 74.79 28.4535 ;
 END
 END vss.gds2462
 PIN vss.gds2463
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 74.732 28.563 74.788 28.763 ;
 RECT 74.564 28.573 74.62 28.773 ;
 RECT 74.06 28.563 74.116 28.763 ;
 RECT 73.892 28.573 73.948 28.773 ;
 RECT 73.388 28.563 73.444 28.763 ;
 RECT 73.22 28.573 73.276 28.773 ;
 RECT 72.716 28.563 72.772 28.763 ;
 RECT 72.548 28.573 72.604 28.773 ;
 RECT 72.044 28.563 72.1 28.763 ;
 RECT 71.876 28.573 71.932 28.773 ;
 RECT 71.372 28.563 71.428 28.763 ;
 RECT 71.204 28.573 71.26 28.773 ;
 RECT 70.7 28.563 70.756 28.763 ;
 RECT 70.532 28.573 70.588 28.773 ;
 RECT 74.396 25.801 74.452 26.001 ;
 RECT 74.228 25.801 74.284 26.001 ;
 RECT 74.564 25.816 74.62 26.016 ;
 RECT 74.732 25.816 74.788 26.016 ;
 RECT 73.724 25.801 73.78 26.001 ;
 RECT 73.556 25.801 73.612 26.001 ;
 RECT 73.892 25.816 73.948 26.016 ;
 RECT 74.06 25.816 74.116 26.016 ;
 RECT 73.052 25.801 73.108 26.001 ;
 RECT 72.884 25.801 72.94 26.001 ;
 RECT 73.22 25.816 73.276 26.016 ;
 RECT 73.388 25.816 73.444 26.016 ;
 RECT 72.38 25.801 72.436 26.001 ;
 RECT 72.212 25.801 72.268 26.001 ;
 RECT 72.548 25.816 72.604 26.016 ;
 RECT 72.716 25.816 72.772 26.016 ;
 RECT 71.708 25.801 71.764 26.001 ;
 RECT 71.54 25.801 71.596 26.001 ;
 RECT 71.876 25.816 71.932 26.016 ;
 RECT 72.044 25.816 72.1 26.016 ;
 RECT 71.036 25.801 71.092 26.001 ;
 RECT 70.868 25.801 70.924 26.001 ;
 RECT 71.204 25.816 71.26 26.016 ;
 RECT 71.372 25.816 71.428 26.016 ;
 RECT 70.364 25.801 70.42 26.001 ;
 RECT 70.532 25.816 70.588 26.016 ;
 RECT 70.7 25.816 70.756 26.016 ;
 RECT 74.396 26.875 74.452 27.075 ;
 RECT 74.228 26.875 74.284 27.075 ;
 RECT 74.564 26.875 74.62 27.075 ;
 RECT 73.724 26.875 73.78 27.075 ;
 RECT 73.556 26.875 73.612 27.075 ;
 RECT 74.06 26.875 74.116 27.075 ;
 RECT 73.892 26.875 73.948 27.075 ;
 RECT 73.052 26.875 73.108 27.075 ;
 RECT 72.884 26.875 72.94 27.075 ;
 RECT 73.388 26.875 73.444 27.075 ;
 RECT 73.22 26.875 73.276 27.075 ;
 RECT 72.38 26.875 72.436 27.075 ;
 RECT 72.212 26.875 72.268 27.075 ;
 RECT 72.716 26.875 72.772 27.075 ;
 RECT 72.548 26.875 72.604 27.075 ;
 RECT 71.708 26.875 71.764 27.075 ;
 RECT 71.54 26.875 71.596 27.075 ;
 RECT 72.044 26.875 72.1 27.075 ;
 RECT 71.876 26.875 71.932 27.075 ;
 RECT 71.036 26.875 71.092 27.075 ;
 RECT 70.868 26.875 70.924 27.075 ;
 RECT 71.372 26.875 71.428 27.075 ;
 RECT 71.204 26.875 71.26 27.075 ;
 RECT 70.364 26.875 70.42 27.075 ;
 RECT 70.7 26.875 70.756 27.075 ;
 RECT 70.532 26.875 70.588 27.075 ;
 RECT 74.732 26.875 74.788 27.075 ;
 END
 END vss.gds2463
 PIN vss.gds2464
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 32.917 2.962 33.117 ;
 END
 END vss.gds2464
 PIN vss.gds2465
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 35.437 2.962 35.637 ;
 END
 END vss.gds2465
 PIN vss.gds2466
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 35.036 3.142 35.236 ;
 END
 END vss.gds2466
 PIN vss.gds2467
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 33.776 3.142 33.976 ;
 END
 END vss.gds2467
 PIN vss.gds2468
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 31.256 3.142 31.456 ;
 END
 END vss.gds2468
 PIN vss.gds2469
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 32.516 3.142 32.716 ;
 END
 END vss.gds2469
 PIN vss.gds2470
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 34.177 2.962 34.377 ;
 END
 END vss.gds2470
 PIN vss.gds2471
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.442 30.621 4.482 30.821 ;
 END
 END vss.gds2471
 PIN vss.gds2472
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 31.657 2.962 31.857 ;
 END
 END vss.gds2472
 PIN vss.gds2473
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.286 31.027 3.326 31.227 ;
 END
 END vss.gds2473
 PIN vss.gds2474
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.754 33.547 3.794 33.747 ;
 END
 END vss.gds2474
 PIN vss.gds2475
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.57 30.824 4.61 31.024 ;
 END
 END vss.gds2475
 PIN vss.gds2476
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.414 31.303 3.454 31.503 ;
 END
 END vss.gds2476
 PIN vss.gds2477
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 33.547 5.074 33.747 ;
 END
 END vss.gds2477
 PIN vss.gds2478
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.562 30.7245 3.602 30.9245 ;
 END
 END vss.gds2478
 PIN vss.gds2479
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 33.141 0.942 33.341 ;
 END
 END vss.gds2479
 PIN vss.gds2480
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 33.547 4.194 33.747 ;
 END
 END vss.gds2480
 PIN vss.gds2481
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 33.2415 0.718 33.4415 ;
 END
 END vss.gds2481
 PIN vss.gds2482
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 33.342 0.602 33.542 ;
 END
 END vss.gds2482
 PIN vss.gds2483
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 33.3755 2.122 33.5755 ;
 END
 END vss.gds2483
 PIN vss.gds2484
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 33.685 1.282 33.885 ;
 END
 END vss.gds2484
 PIN vss.gds2485
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 33.2895 1.462 33.4895 ;
 END
 END vss.gds2485
 PIN vss.gds2486
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 32.852 2.302 33.052 ;
 END
 END vss.gds2486
 PIN vss.gds2487
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 33.4435 4.002 33.6435 ;
 END
 END vss.gds2487
 PIN vss.gds2488
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 33.4435 5.282 33.6435 ;
 END
 END vss.gds2488
 PIN vss.gds2489
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 33.5315 0.29 33.7315 ;
 END
 END vss.gds2489
 PIN vss.gds2490
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 3.332 30.489 3.388 30.689 ;
 RECT 2.408 31.6575 2.464 31.8575 ;
 RECT 2.576 31.6575 2.632 31.8575 ;
 RECT 2.996 31.6575 3.052 31.8575 ;
 RECT 3.332 31.749 3.388 31.949 ;
 RECT 3.5 31.7055 3.556 31.9055 ;
 RECT 0.98 31.5725 1.036 31.7725 ;
 RECT 2.072 31.573 2.128 31.773 ;
 RECT 2.576 32.9175 2.632 33.1175 ;
 RECT 2.408 32.9175 2.464 33.1175 ;
 RECT 2.996 32.9175 3.052 33.1175 ;
 RECT 3.332 33.009 3.388 33.209 ;
 RECT 2.408 34.1775 2.464 34.3775 ;
 RECT 2.576 34.1775 2.632 34.3775 ;
 RECT 2.996 34.1775 3.052 34.3775 ;
 RECT 3.332 34.269 3.388 34.469 ;
 RECT 3.5 34.2255 3.556 34.4255 ;
 RECT 0.98 34.0925 1.036 34.2925 ;
 RECT 2.072 34.093 2.128 34.293 ;
 RECT 2.576 35.4375 2.632 35.6375 ;
 RECT 2.408 35.4375 2.464 35.6375 ;
 RECT 2.996 35.4375 3.052 35.6375 ;
 RECT 0.812 30.489 0.868 30.689 ;
 RECT 0.812 33.009 0.868 33.209 ;
 RECT 0.98 35.3525 1.036 35.5525 ;
 RECT 2.072 35.353 2.128 35.553 ;
 RECT 0.392 35.443 0.448 35.643 ;
 RECT 0.644 35.443 0.7 35.643 ;
 RECT 1.232 35.443 1.288 35.643 ;
 RECT 1.4 35.443 1.456 35.643 ;
 RECT 1.568 35.443 1.624 35.643 ;
 RECT 1.82 35.443 1.876 35.643 ;
 RECT 2.24 35.443 2.296 35.643 ;
 RECT 2.744 35.353 2.8 35.553 ;
 RECT 3.164 35.443 3.22 35.643 ;
 RECT 3.5 32.9655 3.556 33.1655 ;
 RECT 0.392 32.923 0.448 33.123 ;
 RECT 0.644 32.923 0.7 33.123 ;
 RECT 1.232 32.923 1.288 33.123 ;
 RECT 0.98 32.8325 1.036 33.0325 ;
 RECT 1.4 32.923 1.456 33.123 ;
 RECT 1.568 32.923 1.624 33.123 ;
 RECT 2.072 32.833 2.128 33.033 ;
 RECT 1.82 32.923 1.876 33.123 ;
 RECT 2.744 32.833 2.8 33.033 ;
 RECT 3.164 32.923 3.22 33.123 ;
 RECT 2.24 32.923 2.296 33.123 ;
 RECT 3.92 35.443 3.976 35.643 ;
 RECT 0.392 34.183 0.448 34.383 ;
 RECT 0.812 34.269 0.868 34.469 ;
 RECT 0.644 34.183 0.7 34.383 ;
 RECT 1.232 34.183 1.288 34.383 ;
 RECT 1.4 34.183 1.456 34.383 ;
 RECT 1.568 34.183 1.624 34.383 ;
 RECT 1.82 34.183 1.876 34.383 ;
 RECT 2.24 34.183 2.296 34.383 ;
 RECT 2.744 34.093 2.8 34.293 ;
 RECT 3.164 34.183 3.22 34.383 ;
 RECT 3.92 34.183 3.976 34.383 ;
 RECT 3.752 34.453 3.808 34.653 ;
 RECT 4.508 34.3825 4.564 34.5825 ;
 RECT 3.92 32.923 3.976 33.123 ;
 RECT 3.752 33.193 3.808 33.393 ;
 RECT 4.508 33.1225 4.564 33.3225 ;
 RECT 0.392 31.663 0.448 31.863 ;
 RECT 0.812 31.749 0.868 31.949 ;
 RECT 0.644 31.663 0.7 31.863 ;
 RECT 1.232 31.663 1.288 31.863 ;
 RECT 1.4 31.663 1.456 31.863 ;
 RECT 1.568 31.663 1.624 31.863 ;
 RECT 1.82 31.663 1.876 31.863 ;
 RECT 2.24 31.663 2.296 31.863 ;
 RECT 2.744 31.573 2.8 31.773 ;
 RECT 3.164 31.663 3.22 31.863 ;
 RECT 3.92 31.663 3.976 31.863 ;
 RECT 3.752 31.933 3.808 32.133 ;
 RECT 4.508 31.8625 4.564 32.0625 ;
 RECT 3.752 30.673 3.808 30.873 ;
 RECT 4.508 30.6025 4.564 30.8025 ;
 END
 END vss.gds2490
 PIN vss.gds2491
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.134 31.2435 10.194 31.4435 ;
 END
 END vss.gds2491
 PIN vss.gds2492
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.966 31.2435 10.026 31.4435 ;
 END
 END vss.gds2492
 PIN vss.gds2493
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.798 31.2435 9.858 31.4435 ;
 END
 END vss.gds2493
 PIN vss.gds2494
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.462 31.2435 9.522 31.4435 ;
 END
 END vss.gds2494
 PIN vss.gds2495
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.294 31.2435 9.354 31.4435 ;
 END
 END vss.gds2495
 PIN vss.gds2496
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.79 31.2435 8.85 31.4435 ;
 END
 END vss.gds2496
 PIN vss.gds2497
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.622 31.2435 8.682 31.4435 ;
 END
 END vss.gds2497
 PIN vss.gds2498
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.454 31.2435 8.514 31.4435 ;
 END
 END vss.gds2498
 PIN vss.gds2499
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.118 31.2435 8.178 31.4435 ;
 END
 END vss.gds2499
 PIN vss.gds2500
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.95 31.2435 8.01 31.4435 ;
 END
 END vss.gds2500
 PIN vss.gds2501
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.782 31.2435 7.842 31.4435 ;
 END
 END vss.gds2501
 PIN vss.gds2502
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.126 31.2435 9.186 31.4435 ;
 END
 END vss.gds2502
 PIN vss.gds2503
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.446 31.2435 7.506 31.4435 ;
 END
 END vss.gds2503
 PIN vss.gds2504
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.278 31.2435 7.338 31.4435 ;
 END
 END vss.gds2504
 PIN vss.gds2505
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 33.0075 9.69 33.2075 ;
 END
 END vss.gds2505
 PIN vss.gds2506
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 33.0075 9.018 33.2075 ;
 END
 END vss.gds2506
 PIN vss.gds2507
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.11 31.2435 7.17 31.4435 ;
 END
 END vss.gds2507
 PIN vss.gds2508
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 33.344 6.178 33.544 ;
 END
 END vss.gds2508
 PIN vss.gds2509
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 33.547 5.474 33.747 ;
 END
 END vss.gds2509
 PIN vss.gds2510
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 33.0075 8.346 33.2075 ;
 END
 END vss.gds2510
 PIN vss.gds2511
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 33.0075 7.674 33.2075 ;
 END
 END vss.gds2511
 PIN vss.gds2512
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 33.547 5.73 33.747 ;
 END
 END vss.gds2512
 PIN vss.gds2513
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 33.547 5.986 33.747 ;
 END
 END vss.gds2513
 PIN vss.gds2514
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 33.343 6.434 33.543 ;
 END
 END vss.gds2514
 PIN vss.gds2515
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 6.524 35.436 6.58 35.636 ;
 RECT 6.608 34.453 6.664 34.653 ;
 RECT 6.524 34.176 6.58 34.376 ;
 RECT 6.692 34.326 6.748 34.526 ;
 RECT 6.692 33.066 6.748 33.266 ;
 RECT 6.524 32.916 6.58 33.116 ;
 RECT 6.608 33.193 6.664 33.393 ;
 RECT 6.608 31.933 6.664 32.133 ;
 RECT 6.524 31.656 6.58 31.856 ;
 RECT 6.692 31.806 6.748 32.006 ;
 RECT 6.692 30.546 6.748 30.746 ;
 RECT 6.608 30.673 6.664 30.873 ;
 END
 END vss.gds2515
 PIN vss.gds2516
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 32.162 13.898 32.362 ;
 END
 END vss.gds2516
 PIN vss.gds2517
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 32.202 14.87 32.402 ;
 END
 END vss.gds2517
 PIN vss.gds2518
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 33.422 13.898 33.622 ;
 END
 END vss.gds2518
 PIN vss.gds2519
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 33.462 14.87 33.662 ;
 END
 END vss.gds2519
 PIN vss.gds2520
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 34.682 13.898 34.882 ;
 END
 END vss.gds2520
 PIN vss.gds2521
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 34.722 14.87 34.922 ;
 END
 END vss.gds2521
 PIN vss.gds2522
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 30.902 13.898 31.102 ;
 END
 END vss.gds2522
 PIN vss.gds2523
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 30.942 14.87 31.142 ;
 END
 END vss.gds2523
 PIN vss.gds2524
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.15 31.2435 12.21 31.4435 ;
 END
 END vss.gds2524
 PIN vss.gds2525
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.982 31.2435 12.042 31.4435 ;
 END
 END vss.gds2525
 PIN vss.gds2526
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.814 31.2435 11.874 31.4435 ;
 END
 END vss.gds2526
 PIN vss.gds2527
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.478 31.2435 11.538 31.4435 ;
 END
 END vss.gds2527
 PIN vss.gds2528
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.31 31.2435 11.37 31.4435 ;
 END
 END vss.gds2528
 PIN vss.gds2529
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.142 31.2435 11.202 31.4435 ;
 END
 END vss.gds2529
 PIN vss.gds2530
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.806 31.2435 10.866 31.4435 ;
 END
 END vss.gds2530
 PIN vss.gds2531
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.638 31.2435 10.698 31.4435 ;
 END
 END vss.gds2531
 PIN vss.gds2532
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.47 31.2435 10.53 31.4435 ;
 END
 END vss.gds2532
 PIN vss.gds2533
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 31.9295 13.058 32.1295 ;
 END
 END vss.gds2533
 PIN vss.gds2534
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.262 34.236 13.318 34.436 ;
 END
 END vss.gds2534
 PIN vss.gds2535
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 33.0075 11.706 33.2075 ;
 END
 END vss.gds2535
 PIN vss.gds2536
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 33.0075 11.034 33.2075 ;
 END
 END vss.gds2536
 PIN vss.gds2537
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 33.0075 10.362 33.2075 ;
 END
 END vss.gds2537
 PIN vss.gds2538
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 33.173 15.162 33.373 ;
 END
 END vss.gds2538
 PIN vss.gds2539
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 33.173 14.498 33.373 ;
 END
 END vss.gds2539
 PIN vss.gds2540
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 33.0075 13.658 33.2075 ;
 END
 END vss.gds2540
 PIN vss.gds2541
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 32.845 12.378 33.045 ;
 END
 END vss.gds2541
 PIN vss.gds2542
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 33.547 12.59 33.747 ;
 END
 END vss.gds2542
 PIN vss.gds2543
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 33.1635 12.818 33.3635 ;
 END
 END vss.gds2543
 PIN vss.gds2544
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 14 31.08 14.056 31.253 ;
 RECT 14.168 31.053 14.224 31.253 ;
 RECT 14 32.34 14.056 32.513 ;
 RECT 14.168 32.313 14.224 32.513 ;
 RECT 14 33.6 14.056 33.773 ;
 RECT 14.168 33.573 14.224 33.773 ;
 RECT 14 34.86 14.056 35.033 ;
 RECT 14.168 34.833 14.224 35.033 ;
 RECT 14.336 31.673 14.392 31.873 ;
 RECT 14.168 31.673 14.224 31.873 ;
 RECT 14.336 32.933 14.392 33.133 ;
 RECT 14.168 32.933 14.224 33.133 ;
 RECT 14.336 34.193 14.392 34.393 ;
 RECT 14.168 34.193 14.224 34.393 ;
 RECT 15.008 34.403 15.064 34.603 ;
 RECT 14.84 34.877 14.896 35.042 ;
 RECT 14.672 34.877 14.728 35.042 ;
 RECT 13.664 34.327 13.72 34.527 ;
 RECT 13.664 33.067 13.72 33.267 ;
 RECT 15.008 33.143 15.064 33.343 ;
 RECT 14.84 33.617 14.896 33.782 ;
 RECT 14.672 33.617 14.728 33.782 ;
 RECT 13.664 31.807 13.72 32.007 ;
 RECT 15.008 31.883 15.064 32.083 ;
 RECT 14.84 32.357 14.896 32.522 ;
 RECT 14.672 32.357 14.728 32.522 ;
 RECT 13.664 30.547 13.72 30.747 ;
 RECT 15.008 30.623 15.064 30.823 ;
 RECT 14.84 31.097 14.896 31.262 ;
 RECT 14.672 31.097 14.728 31.262 ;
 RECT 15.176 31.3235 15.232 31.5235 ;
 RECT 12.824 31.108 12.88 31.308 ;
 RECT 13.496 31.119 13.552 31.319 ;
 RECT 13.328 31.057 13.384 31.257 ;
 RECT 13.16 31.108 13.216 31.308 ;
 RECT 12.488 31.138 12.544 31.338 ;
 RECT 12.992 31.108 13.048 31.308 ;
 RECT 12.656 31.138 12.712 31.338 ;
 END
 END vss.gds2544
 PIN vss.gds2545
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 34.92 15.418 35.12 ;
 END
 END vss.gds2545
 PIN vss.gds2546
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.438 33.8195 17.494 34.0195 ;
 END
 END vss.gds2546
 PIN vss.gds2547
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 33.0075 20.274 33.2075 ;
 END
 END vss.gds2547
 PIN vss.gds2548
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.702 31.2435 18.762 31.4435 ;
 END
 END vss.gds2548
 PIN vss.gds2549
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.038 31.2435 19.098 31.4435 ;
 END
 END vss.gds2549
 PIN vss.gds2550
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.206 31.2435 19.266 31.4435 ;
 END
 END vss.gds2550
 PIN vss.gds2551
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.374 31.2435 19.434 31.4435 ;
 END
 END vss.gds2551
 PIN vss.gds2552
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.71 31.2435 19.77 31.4435 ;
 END
 END vss.gds2552
 PIN vss.gds2553
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.878 31.2435 19.938 31.4435 ;
 END
 END vss.gds2553
 PIN vss.gds2554
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.534 31.2435 18.594 31.4435 ;
 END
 END vss.gds2554
 PIN vss.gds2555
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 31.716 16.814 31.916 ;
 END
 END vss.gds2555
 PIN vss.gds2556
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 34.177 16.146 34.377 ;
 END
 END vss.gds2556
 PIN vss.gds2557
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 35.437 16.146 35.637 ;
 END
 END vss.gds2557
 PIN vss.gds2558
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 32.917 16.146 33.117 ;
 END
 END vss.gds2558
 PIN vss.gds2559
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 31.657 16.146 31.857 ;
 END
 END vss.gds2559
 PIN vss.gds2560
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.366 31.2435 18.426 31.4435 ;
 END
 END vss.gds2560
 PIN vss.gds2561
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 34.9275 17.314 35.1275 ;
 END
 END vss.gds2561
 PIN vss.gds2562
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.986 31.027 18.026 31.227 ;
 END
 END vss.gds2562
 PIN vss.gds2563
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 33.0075 18.93 33.2075 ;
 END
 END vss.gds2563
 PIN vss.gds2564
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 33.0075 19.602 33.2075 ;
 END
 END vss.gds2564
 PIN vss.gds2565
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 32.9665 16.994 33.1665 ;
 END
 END vss.gds2565
 PIN vss.gds2566
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.046 31.2435 20.106 31.4435 ;
 END
 END vss.gds2566
 PIN vss.gds2567
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 33.173 15.842 33.373 ;
 END
 END vss.gds2567
 PIN vss.gds2568
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 32.845 18.258 33.045 ;
 END
 END vss.gds2568
 PIN vss.gds2569
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 33.1635 17.834 33.3635 ;
 END
 END vss.gds2569
 PIN vss.gds2570
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 33.3755 16.49 33.5755 ;
 END
 END vss.gds2570
 PIN vss.gds2571
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 16.52 31.1 16.576 31.253 ;
 RECT 15.764 31.097 15.82 31.262 ;
 RECT 15.596 31.097 15.652 31.262 ;
 RECT 15.596 31.324 15.652 31.524 ;
 RECT 15.848 31.327 15.904 31.527 ;
 RECT 16.52 32.36 16.576 32.513 ;
 RECT 15.764 32.357 15.82 32.522 ;
 RECT 15.596 32.357 15.652 32.522 ;
 RECT 15.596 32.584 15.652 32.784 ;
 RECT 15.848 32.587 15.904 32.787 ;
 RECT 16.52 33.62 16.576 33.773 ;
 RECT 15.764 33.617 15.82 33.782 ;
 RECT 15.596 33.617 15.652 33.782 ;
 RECT 15.596 33.844 15.652 34.044 ;
 RECT 15.848 33.847 15.904 34.047 ;
 RECT 16.52 34.88 16.576 35.033 ;
 RECT 15.764 34.877 15.82 35.042 ;
 RECT 15.596 34.877 15.652 35.042 ;
 RECT 15.596 35.104 15.652 35.304 ;
 RECT 15.848 35.107 15.904 35.307 ;
 RECT 15.428 34.403 15.484 34.603 ;
 RECT 16.352 34.5035 16.408 34.7035 ;
 RECT 16.856 34.2515 16.912 34.4515 ;
 RECT 16.352 33.2435 16.408 33.4435 ;
 RECT 16.856 32.9915 16.912 33.1915 ;
 RECT 16.352 31.9835 16.408 32.1835 ;
 RECT 16.856 31.7315 16.912 31.9315 ;
 RECT 16.856 30.4715 16.912 30.6715 ;
 RECT 16.352 30.7235 16.408 30.9235 ;
 RECT 15.428 33.143 15.484 33.343 ;
 RECT 15.428 31.883 15.484 32.083 ;
 RECT 15.428 30.623 15.484 30.823 ;
 RECT 17.864 31.138 17.92 31.338 ;
 RECT 17.696 31.1455 17.752 31.3455 ;
 RECT 17.528 31.138 17.584 31.338 ;
 RECT 17.36 31.138 17.416 31.338 ;
 RECT 17.192 31.138 17.248 31.338 ;
 RECT 18.032 31.138 18.088 31.338 ;
 RECT 17.024 31.253 17.08 31.453 ;
 END
 END vss.gds2571
 PIN vss.gds2572
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.17 31.2435 25.23 31.4435 ;
 END
 END vss.gds2572
 PIN vss.gds2573
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.002 31.2435 25.062 31.4435 ;
 END
 END vss.gds2573
 PIN vss.gds2574
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.834 31.2435 24.894 31.4435 ;
 END
 END vss.gds2574
 PIN vss.gds2575
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.498 31.2435 24.558 31.4435 ;
 END
 END vss.gds2575
 PIN vss.gds2576
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.33 31.2435 24.39 31.4435 ;
 END
 END vss.gds2576
 PIN vss.gds2577
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.162 31.2435 24.222 31.4435 ;
 END
 END vss.gds2577
 PIN vss.gds2578
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.382 31.2435 20.442 31.4435 ;
 END
 END vss.gds2578
 PIN vss.gds2579
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.55 31.2435 20.61 31.4435 ;
 END
 END vss.gds2579
 PIN vss.gds2580
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.718 31.2435 20.778 31.4435 ;
 END
 END vss.gds2580
 PIN vss.gds2581
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.054 31.2435 21.114 31.4435 ;
 END
 END vss.gds2581
 PIN vss.gds2582
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.222 31.2435 21.282 31.4435 ;
 END
 END vss.gds2582
 PIN vss.gds2583
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.39 31.2435 21.45 31.4435 ;
 END
 END vss.gds2583
 PIN vss.gds2584
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.726 31.2435 21.786 31.4435 ;
 END
 END vss.gds2584
 PIN vss.gds2585
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.894 31.2435 21.954 31.4435 ;
 END
 END vss.gds2585
 PIN vss.gds2586
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.062 31.2435 22.122 31.4435 ;
 END
 END vss.gds2586
 PIN vss.gds2587
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 33.0075 24.726 33.2075 ;
 END
 END vss.gds2587
 PIN vss.gds2588
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 33.0075 21.618 33.2075 ;
 END
 END vss.gds2588
 PIN vss.gds2589
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 33.0075 20.946 33.2075 ;
 END
 END vss.gds2589
 PIN vss.gds2590
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 33.0075 22.29 33.2075 ;
 END
 END vss.gds2590
 PIN vss.gds2591
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.398 31.2435 22.458 31.4435 ;
 END
 END vss.gds2591
 PIN vss.gds2592
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.566 31.2435 22.626 31.4435 ;
 END
 END vss.gds2592
 PIN vss.gds2593
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.734 31.2435 22.794 31.4435 ;
 END
 END vss.gds2593
 PIN vss.gds2594
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.07 31.2435 23.13 31.4435 ;
 END
 END vss.gds2594
 PIN vss.gds2595
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.238 31.2435 23.298 31.4435 ;
 END
 END vss.gds2595
 PIN vss.gds2596
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.406 31.2435 23.466 31.4435 ;
 END
 END vss.gds2596
 PIN vss.gds2597
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 33.0075 22.962 33.2075 ;
 END
 END vss.gds2597
 PIN vss.gds2598
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 33.0075 23.634 33.2075 ;
 END
 END vss.gds2598
 PIN vss.gds2599
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 23.912 34.34 23.968 34.54 ;
 RECT 23.912 33.08 23.968 33.28 ;
 RECT 23.912 31.82 23.968 32.02 ;
 RECT 23.912 30.56 23.968 30.76 ;
 RECT 23.744 33.08 23.8 33.28 ;
 END
 END vss.gds2599
 PIN vss.gds2600
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.202 31.2435 29.262 31.4435 ;
 END
 END vss.gds2600
 PIN vss.gds2601
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.034 31.2435 29.094 31.4435 ;
 END
 END vss.gds2601
 PIN vss.gds2602
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.866 31.2435 28.926 31.4435 ;
 END
 END vss.gds2602
 PIN vss.gds2603
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.53 31.2435 28.59 31.4435 ;
 END
 END vss.gds2603
 PIN vss.gds2604
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.362 31.2435 28.422 31.4435 ;
 END
 END vss.gds2604
 PIN vss.gds2605
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.194 31.2435 28.254 31.4435 ;
 END
 END vss.gds2605
 PIN vss.gds2606
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.858 31.2435 27.918 31.4435 ;
 END
 END vss.gds2606
 PIN vss.gds2607
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.69 31.2435 27.75 31.4435 ;
 END
 END vss.gds2607
 PIN vss.gds2608
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.522 31.2435 27.582 31.4435 ;
 END
 END vss.gds2608
 PIN vss.gds2609
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.186 31.2435 27.246 31.4435 ;
 END
 END vss.gds2609
 PIN vss.gds2610
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.018 31.2435 27.078 31.4435 ;
 END
 END vss.gds2610
 PIN vss.gds2611
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.85 31.2435 26.91 31.4435 ;
 END
 END vss.gds2611
 PIN vss.gds2612
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.514 31.2435 26.574 31.4435 ;
 END
 END vss.gds2612
 PIN vss.gds2613
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.346 31.2435 26.406 31.4435 ;
 END
 END vss.gds2613
 PIN vss.gds2614
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.178 31.2435 26.238 31.4435 ;
 END
 END vss.gds2614
 PIN vss.gds2615
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.842 31.2435 25.902 31.4435 ;
 END
 END vss.gds2615
 PIN vss.gds2616
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.674 31.2435 25.734 31.4435 ;
 END
 END vss.gds2616
 PIN vss.gds2617
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.506 31.2435 25.566 31.4435 ;
 END
 END vss.gds2617
 PIN vss.gds2618
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 33.0075 28.758 33.2075 ;
 END
 END vss.gds2618
 PIN vss.gds2619
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 33.0075 28.086 33.2075 ;
 END
 END vss.gds2619
 PIN vss.gds2620
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 33.0075 27.414 33.2075 ;
 END
 END vss.gds2620
 PIN vss.gds2621
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 33.0075 26.742 33.2075 ;
 END
 END vss.gds2621
 PIN vss.gds2622
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 33.0075 26.07 33.2075 ;
 END
 END vss.gds2622
 PIN vss.gds2623
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 33.0075 25.398 33.2075 ;
 END
 END vss.gds2623
 PIN vss.gds2624
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 32.845 29.43 33.045 ;
 END
 END vss.gds2624
 PIN vss.gds2625
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 31.9295 30.11 32.1295 ;
 END
 END vss.gds2625
 PIN vss.gds2626
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 33.1635 29.87 33.3635 ;
 END
 END vss.gds2626
 PIN vss.gds2627
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 33.547 29.642 33.747 ;
 END
 END vss.gds2627
 PIN vss.gds2628
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.876 31.108 29.932 31.308 ;
 RECT 29.708 31.138 29.764 31.338 ;
 RECT 30.212 31.108 30.268 31.308 ;
 RECT 29.54 31.138 29.596 31.338 ;
 RECT 30.044 31.108 30.1 31.308 ;
 END
 END vss.gds2628
 PIN vss.gds2629
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 32.202 31.922 32.402 ;
 END
 END vss.gds2629
 PIN vss.gds2630
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 33.422 30.95 33.622 ;
 END
 END vss.gds2630
 PIN vss.gds2631
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 33.462 31.922 33.662 ;
 END
 END vss.gds2631
 PIN vss.gds2632
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 34.682 30.95 34.882 ;
 END
 END vss.gds2632
 PIN vss.gds2633
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 34.722 31.922 34.922 ;
 END
 END vss.gds2633
 PIN vss.gds2634
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 30.902 30.95 31.102 ;
 END
 END vss.gds2634
 PIN vss.gds2635
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 30.942 31.922 31.142 ;
 END
 END vss.gds2635
 PIN vss.gds2636
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 32.162 30.95 32.362 ;
 END
 END vss.gds2636
 PIN vss.gds2637
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.314 34.236 30.37 34.436 ;
 END
 END vss.gds2637
 PIN vss.gds2638
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.49 33.8195 34.546 34.0195 ;
 END
 END vss.gds2638
 PIN vss.gds2639
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 35.437 33.198 35.637 ;
 END
 END vss.gds2639
 PIN vss.gds2640
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 34.177 33.198 34.377 ;
 END
 END vss.gds2640
 PIN vss.gds2641
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 32.917 33.198 33.117 ;
 END
 END vss.gds2641
 PIN vss.gds2642
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 31.657 33.198 31.857 ;
 END
 END vss.gds2642
 PIN vss.gds2643
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 31.716 33.866 31.916 ;
 END
 END vss.gds2643
 PIN vss.gds2644
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 33.173 32.214 33.373 ;
 END
 END vss.gds2644
 PIN vss.gds2645
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 32.9665 34.046 33.1665 ;
 END
 END vss.gds2645
 PIN vss.gds2646
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 34.9275 34.366 35.1275 ;
 END
 END vss.gds2646
 PIN vss.gds2647
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 34.92 32.47 35.12 ;
 END
 END vss.gds2647
 PIN vss.gds2648
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.038 31.027 35.078 31.227 ;
 END
 END vss.gds2648
 PIN vss.gds2649
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 33.0075 30.71 33.2075 ;
 END
 END vss.gds2649
 PIN vss.gds2650
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 33.173 32.894 33.373 ;
 END
 END vss.gds2650
 PIN vss.gds2651
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 33.3755 33.542 33.5755 ;
 END
 END vss.gds2651
 PIN vss.gds2652
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 33.173 31.55 33.373 ;
 END
 END vss.gds2652
 PIN vss.gds2653
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 33.1635 34.886 33.3635 ;
 END
 END vss.gds2653
 PIN vss.gds2654
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 33.572 31.1 33.628 31.253 ;
 RECT 31.052 31.08 31.108 31.253 ;
 RECT 31.22 31.053 31.276 31.253 ;
 RECT 32.816 31.097 32.872 31.262 ;
 RECT 32.648 31.097 32.704 31.262 ;
 RECT 31.892 31.097 31.948 31.262 ;
 RECT 31.724 31.097 31.78 31.262 ;
 RECT 33.572 32.36 33.628 32.513 ;
 RECT 31.052 32.34 31.108 32.513 ;
 RECT 31.22 32.313 31.276 32.513 ;
 RECT 32.816 32.357 32.872 32.522 ;
 RECT 32.648 32.357 32.704 32.522 ;
 RECT 31.892 32.357 31.948 32.522 ;
 RECT 31.724 32.357 31.78 32.522 ;
 RECT 33.572 33.62 33.628 33.773 ;
 RECT 31.052 33.6 31.108 33.773 ;
 RECT 31.22 33.573 31.276 33.773 ;
 RECT 32.816 33.617 32.872 33.782 ;
 RECT 32.648 33.617 32.704 33.782 ;
 RECT 31.892 33.617 31.948 33.782 ;
 RECT 31.724 33.617 31.78 33.782 ;
 RECT 32.648 31.324 32.704 31.524 ;
 RECT 32.9 31.327 32.956 31.527 ;
 RECT 33.572 34.88 33.628 35.033 ;
 RECT 31.052 34.86 31.108 35.033 ;
 RECT 31.22 34.833 31.276 35.033 ;
 RECT 32.816 34.877 32.872 35.042 ;
 RECT 32.648 34.877 32.704 35.042 ;
 RECT 31.892 34.877 31.948 35.042 ;
 RECT 31.724 34.877 31.78 35.042 ;
 RECT 32.648 32.584 32.704 32.784 ;
 RECT 32.9 32.587 32.956 32.787 ;
 RECT 32.648 33.844 32.704 34.044 ;
 RECT 32.9 33.847 32.956 34.047 ;
 RECT 32.648 35.104 32.704 35.304 ;
 RECT 32.9 35.107 32.956 35.307 ;
 RECT 31.388 31.673 31.444 31.873 ;
 RECT 31.22 31.673 31.276 31.873 ;
 RECT 32.06 31.883 32.116 32.083 ;
 RECT 31.388 34.193 31.444 34.393 ;
 RECT 31.22 34.193 31.276 34.393 ;
 RECT 33.404 34.5035 33.46 34.7035 ;
 RECT 33.908 34.2515 33.964 34.4515 ;
 RECT 30.716 31.807 30.772 32.007 ;
 RECT 32.48 31.883 32.536 32.083 ;
 RECT 33.404 33.2435 33.46 33.4435 ;
 RECT 33.908 32.9915 33.964 33.1915 ;
 RECT 31.388 32.933 31.444 33.133 ;
 RECT 31.22 32.933 31.276 33.133 ;
 RECT 33.404 30.7235 33.46 30.9235 ;
 RECT 33.908 30.4715 33.964 30.6715 ;
 RECT 30.716 34.327 30.772 34.527 ;
 RECT 32.06 34.403 32.116 34.603 ;
 RECT 32.48 34.403 32.536 34.603 ;
 RECT 30.716 33.067 30.772 33.267 ;
 RECT 32.06 33.143 32.116 33.343 ;
 RECT 32.48 33.143 32.536 33.343 ;
 RECT 30.716 30.547 30.772 30.747 ;
 RECT 32.06 30.623 32.116 30.823 ;
 RECT 32.48 30.623 32.536 30.823 ;
 RECT 30.548 31.119 30.604 31.319 ;
 RECT 33.404 31.9835 33.46 32.1835 ;
 RECT 33.908 31.7315 33.964 31.9315 ;
 RECT 34.916 31.138 34.972 31.338 ;
 RECT 32.228 31.3235 32.284 31.5235 ;
 RECT 30.38 31.057 30.436 31.257 ;
 RECT 34.748 31.1455 34.804 31.3455 ;
 RECT 34.58 31.138 34.636 31.338 ;
 RECT 34.412 31.138 34.468 31.338 ;
 RECT 34.244 31.138 34.3 31.338 ;
 RECT 34.076 31.253 34.132 31.453 ;
 RECT 35.084 31.138 35.14 31.338 ;
 END
 END vss.gds2654
 PIN vss.gds2655
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.122 31.2435 40.182 31.4435 ;
 END
 END vss.gds2655
 PIN vss.gds2656
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.754 31.2435 35.814 31.4435 ;
 END
 END vss.gds2656
 PIN vss.gds2657
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.09 31.2435 36.15 31.4435 ;
 END
 END vss.gds2657
 PIN vss.gds2658
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.258 31.2435 36.318 31.4435 ;
 END
 END vss.gds2658
 PIN vss.gds2659
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.426 31.2435 36.486 31.4435 ;
 END
 END vss.gds2659
 PIN vss.gds2660
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 33.0075 36.654 33.2075 ;
 END
 END vss.gds2660
 PIN vss.gds2661
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.762 31.2435 36.822 31.4435 ;
 END
 END vss.gds2661
 PIN vss.gds2662
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.93 31.2435 36.99 31.4435 ;
 END
 END vss.gds2662
 PIN vss.gds2663
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.098 31.2435 37.158 31.4435 ;
 END
 END vss.gds2663
 PIN vss.gds2664
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 33.0075 37.326 33.2075 ;
 END
 END vss.gds2664
 PIN vss.gds2665
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.434 31.2435 37.494 31.4435 ;
 END
 END vss.gds2665
 PIN vss.gds2666
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.602 31.2435 37.662 31.4435 ;
 END
 END vss.gds2666
 PIN vss.gds2667
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.77 31.2435 37.83 31.4435 ;
 END
 END vss.gds2667
 PIN vss.gds2668
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 33.0075 37.998 33.2075 ;
 END
 END vss.gds2668
 PIN vss.gds2669
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.106 31.2435 38.166 31.4435 ;
 END
 END vss.gds2669
 PIN vss.gds2670
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.274 31.2435 38.334 31.4435 ;
 END
 END vss.gds2670
 PIN vss.gds2671
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.442 31.2435 38.502 31.4435 ;
 END
 END vss.gds2671
 PIN vss.gds2672
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.778 31.2435 38.838 31.4435 ;
 END
 END vss.gds2672
 PIN vss.gds2673
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.946 31.2435 39.006 31.4435 ;
 END
 END vss.gds2673
 PIN vss.gds2674
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.45 31.2435 39.51 31.4435 ;
 END
 END vss.gds2674
 PIN vss.gds2675
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.618 31.2435 39.678 31.4435 ;
 END
 END vss.gds2675
 PIN vss.gds2676
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.586 31.2435 35.646 31.4435 ;
 END
 END vss.gds2676
 PIN vss.gds2677
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.786 31.2435 39.846 31.4435 ;
 END
 END vss.gds2677
 PIN vss.gds2678
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.114 31.2435 39.174 31.4435 ;
 END
 END vss.gds2678
 PIN vss.gds2679
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.418 31.2435 35.478 31.4435 ;
 END
 END vss.gds2679
 PIN vss.gds2680
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 33.0075 38.67 33.2075 ;
 END
 END vss.gds2680
 PIN vss.gds2681
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 33.0075 35.982 33.2075 ;
 END
 END vss.gds2681
 PIN vss.gds2682
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 33.0075 40.014 33.2075 ;
 END
 END vss.gds2682
 PIN vss.gds2683
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 32.845 35.31 33.045 ;
 END
 END vss.gds2683
 PIN vss.gds2684
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 33.0075 39.342 33.2075 ;
 END
 END vss.gds2684
 PIN vss.gds2685
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 33.0075 45.138 33.2075 ;
 END
 END vss.gds2685
 PIN vss.gds2686
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.91 31.2435 44.97 31.4435 ;
 END
 END vss.gds2686
 PIN vss.gds2687
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.742 31.2435 44.802 31.4435 ;
 END
 END vss.gds2687
 PIN vss.gds2688
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.574 31.2435 44.634 31.4435 ;
 END
 END vss.gds2688
 PIN vss.gds2689
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 33.0075 44.466 33.2075 ;
 END
 END vss.gds2689
 PIN vss.gds2690
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.238 31.2435 44.298 31.4435 ;
 END
 END vss.gds2690
 PIN vss.gds2691
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.07 31.2435 44.13 31.4435 ;
 END
 END vss.gds2691
 PIN vss.gds2692
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.902 31.2435 43.962 31.4435 ;
 END
 END vss.gds2692
 PIN vss.gds2693
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 33.0075 43.794 33.2075 ;
 END
 END vss.gds2693
 PIN vss.gds2694
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.566 31.2435 43.626 31.4435 ;
 END
 END vss.gds2694
 PIN vss.gds2695
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.398 31.2435 43.458 31.4435 ;
 END
 END vss.gds2695
 PIN vss.gds2696
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.23 31.2435 43.29 31.4435 ;
 END
 END vss.gds2696
 PIN vss.gds2697
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 33.0075 43.122 33.2075 ;
 END
 END vss.gds2697
 PIN vss.gds2698
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.894 31.2435 42.954 31.4435 ;
 END
 END vss.gds2698
 PIN vss.gds2699
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.726 31.2435 42.786 31.4435 ;
 END
 END vss.gds2699
 PIN vss.gds2700
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.558 31.2435 42.618 31.4435 ;
 END
 END vss.gds2700
 PIN vss.gds2701
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 33.0075 42.45 33.2075 ;
 END
 END vss.gds2701
 PIN vss.gds2702
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.222 31.2435 42.282 31.4435 ;
 END
 END vss.gds2702
 PIN vss.gds2703
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.054 31.2435 42.114 31.4435 ;
 END
 END vss.gds2703
 PIN vss.gds2704
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.886 31.2435 41.946 31.4435 ;
 END
 END vss.gds2704
 PIN vss.gds2705
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 33.0075 41.778 33.2075 ;
 END
 END vss.gds2705
 PIN vss.gds2706
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.55 31.2435 41.61 31.4435 ;
 END
 END vss.gds2706
 PIN vss.gds2707
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.382 31.2435 41.442 31.4435 ;
 END
 END vss.gds2707
 PIN vss.gds2708
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.214 31.2435 41.274 31.4435 ;
 END
 END vss.gds2708
 PIN vss.gds2709
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.29 31.2435 40.35 31.4435 ;
 END
 END vss.gds2709
 PIN vss.gds2710
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.458 31.2435 40.518 31.4435 ;
 END
 END vss.gds2710
 PIN vss.gds2711
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 33.0075 40.686 33.2075 ;
 END
 END vss.gds2711
 PIN vss.gds2712
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 40.964 34.34 41.02 34.54 ;
 RECT 40.964 31.82 41.02 32.02 ;
 RECT 40.964 30.56 41.02 30.76 ;
 RECT 40.964 33.08 41.02 33.28 ;
 RECT 40.796 33.08 40.852 33.28 ;
 END
 END vss.gds2712
 PIN vss.gds2713
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 32.202 48.974 32.402 ;
 END
 END vss.gds2713
 PIN vss.gds2714
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 33.462 48.974 33.662 ;
 END
 END vss.gds2714
 PIN vss.gds2715
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 34.722 48.974 34.922 ;
 END
 END vss.gds2715
 PIN vss.gds2716
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 30.942 48.974 31.142 ;
 END
 END vss.gds2716
 PIN vss.gds2717
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 32.162 48.002 32.362 ;
 END
 END vss.gds2717
 PIN vss.gds2718
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 33.422 48.002 33.622 ;
 END
 END vss.gds2718
 PIN vss.gds2719
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 34.682 48.002 34.882 ;
 END
 END vss.gds2719
 PIN vss.gds2720
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.366 34.236 47.422 34.436 ;
 END
 END vss.gds2720
 PIN vss.gds2721
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 32.845 46.482 33.045 ;
 END
 END vss.gds2721
 PIN vss.gds2722
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.254 31.2435 46.314 31.4435 ;
 END
 END vss.gds2722
 PIN vss.gds2723
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.086 31.2435 46.146 31.4435 ;
 END
 END vss.gds2723
 PIN vss.gds2724
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.918 31.2435 45.978 31.4435 ;
 END
 END vss.gds2724
 PIN vss.gds2725
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 33.0075 45.81 33.2075 ;
 END
 END vss.gds2725
 PIN vss.gds2726
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.582 31.2435 45.642 31.4435 ;
 END
 END vss.gds2726
 PIN vss.gds2727
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.414 31.2435 45.474 31.4435 ;
 END
 END vss.gds2727
 PIN vss.gds2728
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.246 31.2435 45.306 31.4435 ;
 END
 END vss.gds2728
 PIN vss.gds2729
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 31.9295 47.162 32.1295 ;
 END
 END vss.gds2729
 PIN vss.gds2730
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 34.92 49.522 35.12 ;
 END
 END vss.gds2730
 PIN vss.gds2731
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 35.437 50.25 35.637 ;
 END
 END vss.gds2731
 PIN vss.gds2732
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 34.177 50.25 34.377 ;
 END
 END vss.gds2732
 PIN vss.gds2733
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 32.917 50.25 33.117 ;
 END
 END vss.gds2733
 PIN vss.gds2734
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 33.1635 46.922 33.3635 ;
 END
 END vss.gds2734
 PIN vss.gds2735
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 33.547 46.694 33.747 ;
 END
 END vss.gds2735
 PIN vss.gds2736
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 33.0075 47.762 33.2075 ;
 END
 END vss.gds2736
 PIN vss.gds2737
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 33.173 49.266 33.373 ;
 END
 END vss.gds2737
 PIN vss.gds2738
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 31.657 50.25 31.857 ;
 END
 END vss.gds2738
 PIN vss.gds2739
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 30.902 48.002 31.102 ;
 END
 END vss.gds2739
 PIN vss.gds2740
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 33.173 48.602 33.373 ;
 END
 END vss.gds2740
 PIN vss.gds2741
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 33.173 49.946 33.373 ;
 END
 END vss.gds2741
 PIN vss.gds2742
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 49.7 31.324 49.756 31.524 ;
 RECT 49.952 31.327 50.008 31.527 ;
 RECT 48.104 31.08 48.16 31.253 ;
 RECT 48.272 31.053 48.328 31.253 ;
 RECT 49.868 31.097 49.924 31.262 ;
 RECT 49.7 31.097 49.756 31.262 ;
 RECT 48.944 31.097 49 31.262 ;
 RECT 48.776 31.097 48.832 31.262 ;
 RECT 48.104 32.34 48.16 32.513 ;
 RECT 48.272 32.313 48.328 32.513 ;
 RECT 49.868 32.357 49.924 32.522 ;
 RECT 49.7 32.357 49.756 32.522 ;
 RECT 48.944 32.357 49 32.522 ;
 RECT 48.776 32.357 48.832 32.522 ;
 RECT 48.104 33.6 48.16 33.773 ;
 RECT 48.272 33.573 48.328 33.773 ;
 RECT 49.868 33.617 49.924 33.782 ;
 RECT 49.7 33.617 49.756 33.782 ;
 RECT 48.944 33.617 49 33.782 ;
 RECT 48.776 33.617 48.832 33.782 ;
 RECT 48.104 34.86 48.16 35.033 ;
 RECT 48.272 34.833 48.328 35.033 ;
 RECT 49.868 34.877 49.924 35.042 ;
 RECT 49.7 34.877 49.756 35.042 ;
 RECT 48.944 34.877 49 35.042 ;
 RECT 48.776 34.877 48.832 35.042 ;
 RECT 49.7 35.104 49.756 35.304 ;
 RECT 49.952 35.107 50.008 35.307 ;
 RECT 49.7 33.844 49.756 34.044 ;
 RECT 49.952 33.847 50.008 34.047 ;
 RECT 49.7 32.584 49.756 32.784 ;
 RECT 49.952 32.587 50.008 32.787 ;
 RECT 48.44 32.933 48.496 33.133 ;
 RECT 48.272 32.933 48.328 33.133 ;
 RECT 49.112 34.403 49.168 34.603 ;
 RECT 49.532 34.403 49.588 34.603 ;
 RECT 48.44 34.193 48.496 34.393 ;
 RECT 48.272 34.193 48.328 34.393 ;
 RECT 47.768 34.327 47.824 34.527 ;
 RECT 47.768 33.067 47.824 33.267 ;
 RECT 49.112 33.143 49.168 33.343 ;
 RECT 49.532 33.143 49.588 33.343 ;
 RECT 49.112 30.623 49.168 30.823 ;
 RECT 49.532 30.623 49.588 30.823 ;
 RECT 49.112 31.883 49.168 32.083 ;
 RECT 49.532 31.883 49.588 32.083 ;
 RECT 48.44 31.673 48.496 31.873 ;
 RECT 48.272 31.673 48.328 31.873 ;
 RECT 47.768 31.807 47.824 32.007 ;
 RECT 47.768 30.547 47.824 30.747 ;
 RECT 47.6 31.119 47.656 31.319 ;
 RECT 49.28 31.3235 49.336 31.5235 ;
 RECT 46.928 31.108 46.984 31.308 ;
 RECT 47.432 31.057 47.488 31.257 ;
 RECT 47.264 31.108 47.32 31.308 ;
 RECT 46.592 31.138 46.648 31.338 ;
 RECT 46.76 31.138 46.816 31.338 ;
 RECT 47.096 31.108 47.152 31.308 ;
 END
 END vss.gds2742
 PIN vss.gds2743
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.542 33.8195 51.598 34.0195 ;
 END
 END vss.gds2743
 PIN vss.gds2744
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 31.716 50.918 31.916 ;
 END
 END vss.gds2744
 PIN vss.gds2745
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.638 31.2435 52.698 31.4435 ;
 END
 END vss.gds2745
 PIN vss.gds2746
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.806 31.2435 52.866 31.4435 ;
 END
 END vss.gds2746
 PIN vss.gds2747
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.142 31.2435 53.202 31.4435 ;
 END
 END vss.gds2747
 PIN vss.gds2748
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.31 31.2435 53.37 31.4435 ;
 END
 END vss.gds2748
 PIN vss.gds2749
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.478 31.2435 53.538 31.4435 ;
 END
 END vss.gds2749
 PIN vss.gds2750
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.814 31.2435 53.874 31.4435 ;
 END
 END vss.gds2750
 PIN vss.gds2751
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.982 31.2435 54.042 31.4435 ;
 END
 END vss.gds2751
 PIN vss.gds2752
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.15 31.2435 54.21 31.4435 ;
 END
 END vss.gds2752
 PIN vss.gds2753
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.486 31.2435 54.546 31.4435 ;
 END
 END vss.gds2753
 PIN vss.gds2754
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.654 31.2435 54.714 31.4435 ;
 END
 END vss.gds2754
 PIN vss.gds2755
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.822 31.2435 54.882 31.4435 ;
 END
 END vss.gds2755
 PIN vss.gds2756
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 33.0075 55.05 33.2075 ;
 END
 END vss.gds2756
 PIN vss.gds2757
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.158 31.2435 55.218 31.4435 ;
 END
 END vss.gds2757
 PIN vss.gds2758
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 33.0075 54.378 33.2075 ;
 END
 END vss.gds2758
 PIN vss.gds2759
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 33.0075 53.706 33.2075 ;
 END
 END vss.gds2759
 PIN vss.gds2760
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.47 31.2435 52.53 31.4435 ;
 END
 END vss.gds2760
 PIN vss.gds2761
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 34.9275 51.418 35.1275 ;
 END
 END vss.gds2761
 PIN vss.gds2762
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.09 31.027 52.13 31.227 ;
 END
 END vss.gds2762
 PIN vss.gds2763
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 32.9665 51.098 33.1665 ;
 END
 END vss.gds2763
 PIN vss.gds2764
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 33.0075 53.034 33.2075 ;
 END
 END vss.gds2764
 PIN vss.gds2765
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 33.1635 51.938 33.3635 ;
 END
 END vss.gds2765
 PIN vss.gds2766
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 33.3755 50.594 33.5755 ;
 END
 END vss.gds2766
 PIN vss.gds2767
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 32.845 52.362 33.045 ;
 END
 END vss.gds2767
 PIN vss.gds2768
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 50.624 31.1 50.68 31.253 ;
 RECT 50.624 32.36 50.68 32.513 ;
 RECT 50.624 33.62 50.68 33.773 ;
 RECT 50.624 34.88 50.68 35.033 ;
 RECT 50.96 31.7315 51.016 31.9315 ;
 RECT 50.456 31.9835 50.512 32.1835 ;
 RECT 50.456 30.7235 50.512 30.9235 ;
 RECT 50.96 30.4715 51.016 30.6715 ;
 RECT 50.456 34.5035 50.512 34.7035 ;
 RECT 50.96 34.2515 51.016 34.4515 ;
 RECT 50.456 33.2435 50.512 33.4435 ;
 RECT 50.96 32.9915 51.016 33.1915 ;
 RECT 51.968 31.138 52.024 31.338 ;
 RECT 51.8 31.1455 51.856 31.3455 ;
 RECT 51.632 31.138 51.688 31.338 ;
 RECT 51.464 31.138 51.52 31.338 ;
 RECT 51.296 31.138 51.352 31.338 ;
 RECT 51.128 31.253 51.184 31.453 ;
 RECT 52.136 31.138 52.192 31.338 ;
 END
 END vss.gds2768
 PIN vss.gds2769
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 33.0075 60.174 33.2075 ;
 END
 END vss.gds2769
 PIN vss.gds2770
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.946 31.2435 60.006 31.4435 ;
 END
 END vss.gds2770
 PIN vss.gds2771
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.778 31.2435 59.838 31.4435 ;
 END
 END vss.gds2771
 PIN vss.gds2772
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.61 31.2435 59.67 31.4435 ;
 END
 END vss.gds2772
 PIN vss.gds2773
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 33.0075 59.502 33.2075 ;
 END
 END vss.gds2773
 PIN vss.gds2774
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.274 31.2435 59.334 31.4435 ;
 END
 END vss.gds2774
 PIN vss.gds2775
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.106 31.2435 59.166 31.4435 ;
 END
 END vss.gds2775
 PIN vss.gds2776
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.938 31.2435 58.998 31.4435 ;
 END
 END vss.gds2776
 PIN vss.gds2777
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 33.0075 58.83 33.2075 ;
 END
 END vss.gds2777
 PIN vss.gds2778
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.602 31.2435 58.662 31.4435 ;
 END
 END vss.gds2778
 PIN vss.gds2779
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.434 31.2435 58.494 31.4435 ;
 END
 END vss.gds2779
 PIN vss.gds2780
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.266 31.2435 58.326 31.4435 ;
 END
 END vss.gds2780
 PIN vss.gds2781
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.326 31.2435 55.386 31.4435 ;
 END
 END vss.gds2781
 PIN vss.gds2782
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.494 31.2435 55.554 31.4435 ;
 END
 END vss.gds2782
 PIN vss.gds2783
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.83 31.2435 55.89 31.4435 ;
 END
 END vss.gds2783
 PIN vss.gds2784
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.998 31.2435 56.058 31.4435 ;
 END
 END vss.gds2784
 PIN vss.gds2785
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.166 31.2435 56.226 31.4435 ;
 END
 END vss.gds2785
 PIN vss.gds2786
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.502 31.2435 56.562 31.4435 ;
 END
 END vss.gds2786
 PIN vss.gds2787
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.67 31.2435 56.73 31.4435 ;
 END
 END vss.gds2787
 PIN vss.gds2788
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.838 31.2435 56.898 31.4435 ;
 END
 END vss.gds2788
 PIN vss.gds2789
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.342 31.2435 57.402 31.4435 ;
 END
 END vss.gds2789
 PIN vss.gds2790
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.51 31.2435 57.57 31.4435 ;
 END
 END vss.gds2790
 PIN vss.gds2791
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 33.0075 55.722 33.2075 ;
 END
 END vss.gds2791
 PIN vss.gds2792
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 33.0075 56.394 33.2075 ;
 END
 END vss.gds2792
 PIN vss.gds2793
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.174 31.2435 57.234 31.4435 ;
 END
 END vss.gds2793
 PIN vss.gds2794
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 33.0075 57.738 33.2075 ;
 END
 END vss.gds2794
 PIN vss.gds2795
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 33.0075 57.066 33.2075 ;
 END
 END vss.gds2795
 PIN vss.gds2796
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 58.016 33.08 58.072 33.28 ;
 RECT 58.016 34.34 58.072 34.54 ;
 RECT 58.016 30.56 58.072 30.76 ;
 RECT 58.016 31.82 58.072 32.02 ;
 RECT 57.848 33.08 57.904 33.28 ;
 END
 END vss.gds2796
 PIN vss.gds2797
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 33.422 65.054 33.622 ;
 END
 END vss.gds2797
 PIN vss.gds2798
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 30.902 65.054 31.102 ;
 END
 END vss.gds2798
 PIN vss.gds2799
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 32.162 65.054 32.362 ;
 END
 END vss.gds2799
 PIN vss.gds2800
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 31.9295 64.214 32.1295 ;
 END
 END vss.gds2800
 PIN vss.gds2801
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.418 34.236 64.474 34.436 ;
 END
 END vss.gds2801
 PIN vss.gds2802
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 32.845 63.534 33.045 ;
 END
 END vss.gds2802
 PIN vss.gds2803
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.306 31.2435 63.366 31.4435 ;
 END
 END vss.gds2803
 PIN vss.gds2804
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.138 31.2435 63.198 31.4435 ;
 END
 END vss.gds2804
 PIN vss.gds2805
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.97 31.2435 63.03 31.4435 ;
 END
 END vss.gds2805
 PIN vss.gds2806
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 33.0075 62.862 33.2075 ;
 END
 END vss.gds2806
 PIN vss.gds2807
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.634 31.2435 62.694 31.4435 ;
 END
 END vss.gds2807
 PIN vss.gds2808
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.466 31.2435 62.526 31.4435 ;
 END
 END vss.gds2808
 PIN vss.gds2809
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.298 31.2435 62.358 31.4435 ;
 END
 END vss.gds2809
 PIN vss.gds2810
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 33.0075 62.19 33.2075 ;
 END
 END vss.gds2810
 PIN vss.gds2811
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.962 31.2435 62.022 31.4435 ;
 END
 END vss.gds2811
 PIN vss.gds2812
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.794 31.2435 61.854 31.4435 ;
 END
 END vss.gds2812
 PIN vss.gds2813
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.626 31.2435 61.686 31.4435 ;
 END
 END vss.gds2813
 PIN vss.gds2814
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 33.0075 61.518 33.2075 ;
 END
 END vss.gds2814
 PIN vss.gds2815
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.29 31.2435 61.35 31.4435 ;
 END
 END vss.gds2815
 PIN vss.gds2816
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.122 31.2435 61.182 31.4435 ;
 END
 END vss.gds2816
 PIN vss.gds2817
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.954 31.2435 61.014 31.4435 ;
 END
 END vss.gds2817
 PIN vss.gds2818
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 33.0075 60.846 33.2075 ;
 END
 END vss.gds2818
 PIN vss.gds2819
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.618 31.2435 60.678 31.4435 ;
 END
 END vss.gds2819
 PIN vss.gds2820
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.45 31.2435 60.51 31.4435 ;
 END
 END vss.gds2820
 PIN vss.gds2821
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.282 31.2435 60.342 31.4435 ;
 END
 END vss.gds2821
 PIN vss.gds2822
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 33.1635 63.974 33.3635 ;
 END
 END vss.gds2822
 PIN vss.gds2823
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 33.547 63.746 33.747 ;
 END
 END vss.gds2823
 PIN vss.gds2824
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 34.682 65.054 34.882 ;
 END
 END vss.gds2824
 PIN vss.gds2825
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 33.0075 64.814 33.2075 ;
 END
 END vss.gds2825
 PIN vss.gds2826
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 65.156 31.08 65.212 31.253 ;
 RECT 65.156 32.34 65.212 32.513 ;
 RECT 65.156 33.6 65.212 33.773 ;
 RECT 65.156 34.86 65.212 35.033 ;
 RECT 64.82 34.327 64.876 34.527 ;
 RECT 64.82 30.547 64.876 30.747 ;
 RECT 64.82 31.807 64.876 32.007 ;
 RECT 64.82 33.067 64.876 33.267 ;
 RECT 64.652 31.119 64.708 31.319 ;
 RECT 63.98 31.108 64.036 31.308 ;
 RECT 63.812 31.138 63.868 31.338 ;
 RECT 64.484 31.057 64.54 31.257 ;
 RECT 64.316 31.108 64.372 31.308 ;
 RECT 63.644 31.138 63.7 31.338 ;
 RECT 64.148 31.108 64.204 31.308 ;
 END
 END vss.gds2826
 PIN vss.gds2827
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 32.202 66.026 32.402 ;
 END
 END vss.gds2827
 PIN vss.gds2828
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 33.462 66.026 33.662 ;
 END
 END vss.gds2828
 PIN vss.gds2829
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 34.722 66.026 34.922 ;
 END
 END vss.gds2829
 PIN vss.gds2830
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 30.942 66.026 31.142 ;
 END
 END vss.gds2830
 PIN vss.gds2831
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 35.437 67.302 35.637 ;
 END
 END vss.gds2831
 PIN vss.gds2832
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 34.177 67.302 34.377 ;
 END
 END vss.gds2832
 PIN vss.gds2833
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 34.92 66.574 35.12 ;
 END
 END vss.gds2833
 PIN vss.gds2834
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.594 33.8195 68.65 34.0195 ;
 END
 END vss.gds2834
 PIN vss.gds2835
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 32.9665 68.15 33.1665 ;
 END
 END vss.gds2835
 PIN vss.gds2836
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.858 31.2435 69.918 31.4435 ;
 END
 END vss.gds2836
 PIN vss.gds2837
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.194 31.2435 70.254 31.4435 ;
 END
 END vss.gds2837
 PIN vss.gds2838
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.142 31.027 69.182 31.227 ;
 END
 END vss.gds2838
 PIN vss.gds2839
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 32.917 67.302 33.117 ;
 END
 END vss.gds2839
 PIN vss.gds2840
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 31.716 67.97 31.916 ;
 END
 END vss.gds2840
 PIN vss.gds2841
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 31.657 67.302 31.857 ;
 END
 END vss.gds2841
 PIN vss.gds2842
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.69 31.2435 69.75 31.4435 ;
 END
 END vss.gds2842
 PIN vss.gds2843
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 33.173 66.318 33.373 ;
 END
 END vss.gds2843
 PIN vss.gds2844
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.522 31.2435 69.582 31.4435 ;
 END
 END vss.gds2844
 PIN vss.gds2845
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 34.9275 68.47 35.1275 ;
 END
 END vss.gds2845
 PIN vss.gds2846
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 33.0075 70.086 33.2075 ;
 END
 END vss.gds2846
 PIN vss.gds2847
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 33.173 66.998 33.373 ;
 END
 END vss.gds2847
 PIN vss.gds2848
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 33.173 65.654 33.373 ;
 END
 END vss.gds2848
 PIN vss.gds2849
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 33.3755 67.646 33.5755 ;
 END
 END vss.gds2849
 PIN vss.gds2850
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 33.1635 68.99 33.3635 ;
 END
 END vss.gds2850
 PIN vss.gds2851
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 32.845 69.414 33.045 ;
 END
 END vss.gds2851
 PIN vss.gds2852
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 66.752 32.584 66.808 32.784 ;
 RECT 67.004 32.587 67.06 32.787 ;
 RECT 67.676 31.1 67.732 31.253 ;
 RECT 65.324 31.053 65.38 31.253 ;
 RECT 66.92 31.097 66.976 31.262 ;
 RECT 66.752 31.097 66.808 31.262 ;
 RECT 65.996 31.097 66.052 31.262 ;
 RECT 65.828 31.097 65.884 31.262 ;
 RECT 67.676 32.36 67.732 32.513 ;
 RECT 65.324 32.313 65.38 32.513 ;
 RECT 66.92 32.357 66.976 32.522 ;
 RECT 66.752 32.357 66.808 32.522 ;
 RECT 65.996 32.357 66.052 32.522 ;
 RECT 65.828 32.357 65.884 32.522 ;
 RECT 67.676 33.62 67.732 33.773 ;
 RECT 65.324 33.573 65.38 33.773 ;
 RECT 66.92 33.617 66.976 33.782 ;
 RECT 66.752 33.617 66.808 33.782 ;
 RECT 65.996 33.617 66.052 33.782 ;
 RECT 65.828 33.617 65.884 33.782 ;
 RECT 66.752 33.844 66.808 34.044 ;
 RECT 67.004 33.847 67.06 34.047 ;
 RECT 67.676 34.88 67.732 35.033 ;
 RECT 65.324 34.833 65.38 35.033 ;
 RECT 66.92 34.877 66.976 35.042 ;
 RECT 66.752 34.877 66.808 35.042 ;
 RECT 65.996 34.877 66.052 35.042 ;
 RECT 65.828 34.877 65.884 35.042 ;
 RECT 66.752 31.324 66.808 31.524 ;
 RECT 67.004 31.327 67.06 31.527 ;
 RECT 66.752 35.104 66.808 35.304 ;
 RECT 67.004 35.107 67.06 35.307 ;
 RECT 65.492 34.193 65.548 34.393 ;
 RECT 65.324 34.193 65.38 34.393 ;
 RECT 66.164 34.403 66.22 34.603 ;
 RECT 66.584 34.403 66.64 34.603 ;
 RECT 67.508 34.5035 67.564 34.7035 ;
 RECT 68.012 34.2515 68.068 34.4515 ;
 RECT 66.164 31.883 66.22 32.083 ;
 RECT 65.492 31.673 65.548 31.873 ;
 RECT 65.324 31.673 65.38 31.873 ;
 RECT 66.584 31.883 66.64 32.083 ;
 RECT 66.164 30.623 66.22 30.823 ;
 RECT 67.508 31.9835 67.564 32.1835 ;
 RECT 68.012 31.7315 68.068 31.9315 ;
 RECT 68.012 32.9915 68.068 33.1915 ;
 RECT 67.508 33.2435 67.564 33.4435 ;
 RECT 66.164 33.143 66.22 33.343 ;
 RECT 66.584 33.143 66.64 33.343 ;
 RECT 65.492 32.933 65.548 33.133 ;
 RECT 65.324 32.933 65.38 33.133 ;
 RECT 66.584 30.623 66.64 30.823 ;
 RECT 67.508 30.7235 67.564 30.9235 ;
 RECT 68.012 30.4715 68.068 30.6715 ;
 RECT 66.332 31.3235 66.388 31.5235 ;
 RECT 69.02 31.138 69.076 31.338 ;
 RECT 68.852 31.1455 68.908 31.3455 ;
 RECT 68.684 31.138 68.74 31.338 ;
 RECT 68.516 31.138 68.572 31.338 ;
 RECT 68.348 31.138 68.404 31.338 ;
 RECT 69.188 31.138 69.244 31.338 ;
 RECT 68.18 31.253 68.236 31.453 ;
 END
 END vss.gds2852
 PIN vss.gds2853
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.362 31.2435 70.422 31.4435 ;
 END
 END vss.gds2853
 PIN vss.gds2854
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.53 31.2435 70.59 31.4435 ;
 END
 END vss.gds2854
 PIN vss.gds2855
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.866 31.2435 70.926 31.4435 ;
 END
 END vss.gds2855
 PIN vss.gds2856
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.034 31.2435 71.094 31.4435 ;
 END
 END vss.gds2856
 PIN vss.gds2857
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.202 31.2435 71.262 31.4435 ;
 END
 END vss.gds2857
 PIN vss.gds2858
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 33.0075 71.43 33.2075 ;
 END
 END vss.gds2858
 PIN vss.gds2859
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.538 31.2435 71.598 31.4435 ;
 END
 END vss.gds2859
 PIN vss.gds2860
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.706 31.2435 71.766 31.4435 ;
 END
 END vss.gds2860
 PIN vss.gds2861
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.874 31.2435 71.934 31.4435 ;
 END
 END vss.gds2861
 PIN vss.gds2862
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 33.0075 72.102 33.2075 ;
 END
 END vss.gds2862
 PIN vss.gds2863
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.21 31.2435 72.27 31.4435 ;
 END
 END vss.gds2863
 PIN vss.gds2864
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.378 31.2435 72.438 31.4435 ;
 END
 END vss.gds2864
 PIN vss.gds2865
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.546 31.2435 72.606 31.4435 ;
 END
 END vss.gds2865
 PIN vss.gds2866
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 33.0075 72.774 33.2075 ;
 END
 END vss.gds2866
 PIN vss.gds2867
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.882 31.2435 72.942 31.4435 ;
 END
 END vss.gds2867
 PIN vss.gds2868
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.05 31.2435 73.11 31.4435 ;
 END
 END vss.gds2868
 PIN vss.gds2869
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.554 31.2435 73.614 31.4435 ;
 END
 END vss.gds2869
 PIN vss.gds2870
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.722 31.2435 73.782 31.4435 ;
 END
 END vss.gds2870
 PIN vss.gds2871
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.89 31.2435 73.95 31.4435 ;
 END
 END vss.gds2871
 PIN vss.gds2872
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.394 31.2435 74.454 31.4435 ;
 END
 END vss.gds2872
 PIN vss.gds2873
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.218 31.2435 73.278 31.4435 ;
 END
 END vss.gds2873
 PIN vss.gds2874
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.562 31.2435 74.622 31.4435 ;
 END
 END vss.gds2874
 PIN vss.gds2875
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.226 31.2435 74.286 31.4435 ;
 END
 END vss.gds2875
 PIN vss.gds2876
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 33.0075 70.758 33.2075 ;
 END
 END vss.gds2876
 PIN vss.gds2877
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 33.0075 73.446 33.2075 ;
 END
 END vss.gds2877
 PIN vss.gds2878
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 33.0075 74.118 33.2075 ;
 END
 END vss.gds2878
 PIN vss.gds2879
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 33.0075 74.79 33.2075 ;
 END
 END vss.gds2879
 PIN vss.gds2880
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 37.957 2.962 38.157 ;
 END
 END vss.gds2880
 PIN vss.gds2881
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 39.217 2.962 39.417 ;
 END
 END vss.gds2881
 PIN vss.gds2882
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 36.296 3.142 36.496 ;
 END
 END vss.gds2882
 PIN vss.gds2883
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 36.697 2.962 36.897 ;
 END
 END vss.gds2883
 PIN vss.gds2884
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 37.556 3.142 37.756 ;
 END
 END vss.gds2884
 PIN vss.gds2885
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 38.816 3.142 39.016 ;
 END
 END vss.gds2885
 PIN vss.gds2886
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 40.076 3.142 40.276 ;
 END
 END vss.gds2886
 PIN vss.gds2887
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.442 35.661 4.482 35.861 ;
 END
 END vss.gds2887
 PIN vss.gds2888
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.286 36.067 3.326 36.267 ;
 END
 END vss.gds2888
 PIN vss.gds2889
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.754 38.587 3.794 38.787 ;
 END
 END vss.gds2889
 PIN vss.gds2890
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.57 35.864 4.61 36.064 ;
 END
 END vss.gds2890
 PIN vss.gds2891
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.414 36.343 3.454 36.543 ;
 END
 END vss.gds2891
 PIN vss.gds2892
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 35.661 4.882 35.861 ;
 END
 END vss.gds2892
 PIN vss.gds2893
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 38.587 5.074 38.787 ;
 END
 END vss.gds2893
 PIN vss.gds2894
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.562 36.343 3.602 36.543 ;
 END
 END vss.gds2894
 PIN vss.gds2895
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 38.181 0.942 38.381 ;
 END
 END vss.gds2895
 PIN vss.gds2896
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 38.587 4.194 38.787 ;
 END
 END vss.gds2896
 PIN vss.gds2897
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 38.2815 0.718 38.4815 ;
 END
 END vss.gds2897
 PIN vss.gds2898
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 38.382 0.602 38.582 ;
 END
 END vss.gds2898
 PIN vss.gds2899
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 38.1905 2.122 38.3905 ;
 END
 END vss.gds2899
 PIN vss.gds2900
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 38.725 1.282 38.925 ;
 END
 END vss.gds2900
 PIN vss.gds2901
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 38.3295 1.462 38.5295 ;
 END
 END vss.gds2901
 PIN vss.gds2902
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 37.892 2.302 38.092 ;
 END
 END vss.gds2902
 PIN vss.gds2903
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 38.4835 4.002 38.6835 ;
 END
 END vss.gds2903
 PIN vss.gds2904
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 38.4835 5.282 38.6835 ;
 END
 END vss.gds2904
 PIN vss.gds2905
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 38.491 0.29 38.691 ;
 END
 END vss.gds2905
 PIN vss.gds2906
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 3.332 35.529 3.388 35.729 ;
 RECT 2.408 36.6975 2.464 36.8975 ;
 RECT 2.576 36.6975 2.632 36.8975 ;
 RECT 2.996 36.6975 3.052 36.8975 ;
 RECT 3.332 36.789 3.388 36.989 ;
 RECT 3.5 36.7455 3.556 36.9455 ;
 RECT 0.98 36.6125 1.036 36.8125 ;
 RECT 2.072 36.613 2.128 36.813 ;
 RECT 2.576 37.9575 2.632 38.1575 ;
 RECT 2.408 37.9575 2.464 38.1575 ;
 RECT 2.996 37.9575 3.052 38.1575 ;
 RECT 3.332 38.049 3.388 38.249 ;
 RECT 2.408 39.2175 2.464 39.4175 ;
 RECT 2.576 39.2175 2.632 39.4175 ;
 RECT 2.996 39.2175 3.052 39.4175 ;
 RECT 3.332 39.309 3.388 39.509 ;
 RECT 3.5 39.2655 3.556 39.4655 ;
 RECT 0.98 39.1325 1.036 39.3325 ;
 RECT 2.072 39.133 2.128 39.333 ;
 RECT 3.5 35.4855 3.556 35.6855 ;
 RECT 0.812 38.049 0.868 38.249 ;
 RECT 0.98 40.3925 1.036 40.5925 ;
 RECT 2.072 40.393 2.128 40.593 ;
 RECT 2.744 40.393 2.8 40.593 ;
 RECT 3.5 38.0055 3.556 38.2055 ;
 RECT 0.392 37.963 0.448 38.163 ;
 RECT 0.644 37.963 0.7 38.163 ;
 RECT 1.232 37.963 1.288 38.163 ;
 RECT 0.98 37.8725 1.036 38.0725 ;
 RECT 1.4 37.963 1.456 38.163 ;
 RECT 1.568 37.963 1.624 38.163 ;
 RECT 2.072 37.873 2.128 38.073 ;
 RECT 1.82 37.963 1.876 38.163 ;
 RECT 2.744 37.873 2.8 38.073 ;
 RECT 3.164 37.963 3.22 38.163 ;
 RECT 2.24 37.963 2.296 38.163 ;
 RECT 0.812 35.529 0.868 35.729 ;
 RECT 0.392 39.223 0.448 39.423 ;
 RECT 0.812 39.309 0.868 39.509 ;
 RECT 0.644 39.223 0.7 39.423 ;
 RECT 1.232 39.223 1.288 39.423 ;
 RECT 1.4 39.223 1.456 39.423 ;
 RECT 1.568 39.223 1.624 39.423 ;
 RECT 1.82 39.223 1.876 39.423 ;
 RECT 2.24 39.223 2.296 39.423 ;
 RECT 2.744 39.133 2.8 39.333 ;
 RECT 3.164 39.223 3.22 39.423 ;
 RECT 3.92 39.223 3.976 39.423 ;
 RECT 3.752 39.493 3.808 39.693 ;
 RECT 4.508 39.4225 4.564 39.6225 ;
 RECT 3.92 37.963 3.976 38.163 ;
 RECT 3.752 38.233 3.808 38.433 ;
 RECT 4.508 38.1625 4.564 38.3625 ;
 RECT 0.392 36.703 0.448 36.903 ;
 RECT 0.812 36.789 0.868 36.989 ;
 RECT 0.644 36.703 0.7 36.903 ;
 RECT 1.232 36.703 1.288 36.903 ;
 RECT 1.4 36.703 1.456 36.903 ;
 RECT 1.568 36.703 1.624 36.903 ;
 RECT 1.82 36.703 1.876 36.903 ;
 RECT 2.24 36.703 2.296 36.903 ;
 RECT 2.744 36.613 2.8 36.813 ;
 RECT 3.164 36.703 3.22 36.903 ;
 RECT 3.92 36.703 3.976 36.903 ;
 RECT 3.752 36.973 3.808 37.173 ;
 RECT 4.508 36.9025 4.564 37.1025 ;
 RECT 3.752 35.713 3.808 35.913 ;
 RECT 4.508 35.6425 4.564 35.8425 ;
 END
 END vss.gds2906
 PIN vss.gds2907
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.134 36.2835 10.194 36.4835 ;
 END
 END vss.gds2907
 PIN vss.gds2908
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.966 36.2835 10.026 36.4835 ;
 END
 END vss.gds2908
 PIN vss.gds2909
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.798 36.2835 9.858 36.4835 ;
 END
 END vss.gds2909
 PIN vss.gds2910
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.462 36.2835 9.522 36.4835 ;
 END
 END vss.gds2910
 PIN vss.gds2911
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.294 36.2835 9.354 36.4835 ;
 END
 END vss.gds2911
 PIN vss.gds2912
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.79 36.2835 8.85 36.4835 ;
 END
 END vss.gds2912
 PIN vss.gds2913
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.622 36.2835 8.682 36.4835 ;
 END
 END vss.gds2913
 PIN vss.gds2914
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.454 36.2835 8.514 36.4835 ;
 END
 END vss.gds2914
 PIN vss.gds2915
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.118 36.2835 8.178 36.4835 ;
 END
 END vss.gds2915
 PIN vss.gds2916
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.95 36.2835 8.01 36.4835 ;
 END
 END vss.gds2916
 PIN vss.gds2917
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.782 36.2835 7.842 36.4835 ;
 END
 END vss.gds2917
 PIN vss.gds2918
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.126 36.2835 9.186 36.4835 ;
 END
 END vss.gds2918
 PIN vss.gds2919
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.446 36.2835 7.506 36.4835 ;
 END
 END vss.gds2919
 PIN vss.gds2920
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.278 36.2835 7.338 36.4835 ;
 END
 END vss.gds2920
 PIN vss.gds2921
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 38.0475 9.69 38.2475 ;
 END
 END vss.gds2921
 PIN vss.gds2922
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 38.0475 9.018 38.2475 ;
 END
 END vss.gds2922
 PIN vss.gds2923
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.11 36.2835 7.17 36.4835 ;
 END
 END vss.gds2923
 PIN vss.gds2924
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 38.384 6.178 38.584 ;
 END
 END vss.gds2924
 PIN vss.gds2925
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 38.587 5.474 38.787 ;
 END
 END vss.gds2925
 PIN vss.gds2926
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 38.0475 8.346 38.2475 ;
 END
 END vss.gds2926
 PIN vss.gds2927
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 38.0475 7.674 38.2475 ;
 END
 END vss.gds2927
 PIN vss.gds2928
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 38.587 5.73 38.787 ;
 END
 END vss.gds2928
 PIN vss.gds2929
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 38.587 5.986 38.787 ;
 END
 END vss.gds2929
 PIN vss.gds2930
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 38.383 6.434 38.583 ;
 END
 END vss.gds2930
 PIN vss.gds2931
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 6.608 39.493 6.664 39.693 ;
 RECT 6.524 39.216 6.58 39.416 ;
 RECT 6.692 39.366 6.748 39.566 ;
 RECT 6.692 38.106 6.748 38.306 ;
 RECT 6.524 37.956 6.58 38.156 ;
 RECT 6.608 38.233 6.664 38.433 ;
 RECT 6.608 36.973 6.664 37.173 ;
 RECT 6.524 36.696 6.58 36.896 ;
 RECT 6.692 36.846 6.748 37.046 ;
 RECT 6.692 35.586 6.748 35.786 ;
 RECT 6.608 35.713 6.664 35.913 ;
 END
 END vss.gds2931
 PIN vss.gds2932
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 37.202 13.898 37.402 ;
 END
 END vss.gds2932
 PIN vss.gds2933
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 37.242 14.87 37.442 ;
 END
 END vss.gds2933
 PIN vss.gds2934
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 35.942 13.898 36.142 ;
 END
 END vss.gds2934
 PIN vss.gds2935
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 35.982 14.87 36.182 ;
 END
 END vss.gds2935
 PIN vss.gds2936
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 39.722 13.898 39.922 ;
 END
 END vss.gds2936
 PIN vss.gds2937
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 39.762 14.87 39.962 ;
 END
 END vss.gds2937
 PIN vss.gds2938
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 38.462 13.898 38.662 ;
 END
 END vss.gds2938
 PIN vss.gds2939
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 38.502 14.87 38.702 ;
 END
 END vss.gds2939
 PIN vss.gds2940
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.15 36.2835 12.21 36.4835 ;
 END
 END vss.gds2940
 PIN vss.gds2941
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.982 36.2835 12.042 36.4835 ;
 END
 END vss.gds2941
 PIN vss.gds2942
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.814 36.2835 11.874 36.4835 ;
 END
 END vss.gds2942
 PIN vss.gds2943
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.478 36.2835 11.538 36.4835 ;
 END
 END vss.gds2943
 PIN vss.gds2944
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.31 36.2835 11.37 36.4835 ;
 END
 END vss.gds2944
 PIN vss.gds2945
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.142 36.2835 11.202 36.4835 ;
 END
 END vss.gds2945
 PIN vss.gds2946
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.806 36.2835 10.866 36.4835 ;
 END
 END vss.gds2946
 PIN vss.gds2947
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.638 36.2835 10.698 36.4835 ;
 END
 END vss.gds2947
 PIN vss.gds2948
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.47 36.2835 10.53 36.4835 ;
 END
 END vss.gds2948
 PIN vss.gds2949
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 36.9695 13.058 37.1695 ;
 END
 END vss.gds2949
 PIN vss.gds2950
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.262 39.276 13.318 39.476 ;
 END
 END vss.gds2950
 PIN vss.gds2951
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 38.0475 11.706 38.2475 ;
 END
 END vss.gds2951
 PIN vss.gds2952
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 38.0475 11.034 38.2475 ;
 END
 END vss.gds2952
 PIN vss.gds2953
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 38.0475 10.362 38.2475 ;
 END
 END vss.gds2953
 PIN vss.gds2954
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 38.088 15.162 38.288 ;
 END
 END vss.gds2954
 PIN vss.gds2955
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 38.088 14.498 38.288 ;
 END
 END vss.gds2955
 PIN vss.gds2956
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 38.0475 13.658 38.2475 ;
 END
 END vss.gds2956
 PIN vss.gds2957
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 37.885 12.378 38.085 ;
 END
 END vss.gds2957
 PIN vss.gds2958
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 38.587 12.59 38.787 ;
 END
 END vss.gds2958
 PIN vss.gds2959
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 38.2035 12.818 38.4035 ;
 END
 END vss.gds2959
 PIN vss.gds2960
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 14 36.12 14.056 36.293 ;
 RECT 14.168 36.093 14.224 36.293 ;
 RECT 14 37.38 14.056 37.553 ;
 RECT 14.168 37.353 14.224 37.553 ;
 RECT 14 38.64 14.056 38.813 ;
 RECT 14.168 38.613 14.224 38.813 ;
 RECT 14 39.9 14.056 40.073 ;
 RECT 14.168 39.873 14.224 40.073 ;
 RECT 14.336 36.713 14.392 36.913 ;
 RECT 14.168 36.713 14.224 36.913 ;
 RECT 14.336 35.453 14.392 35.653 ;
 RECT 14.168 35.453 14.224 35.653 ;
 RECT 14.336 39.233 14.392 39.433 ;
 RECT 14.168 39.233 14.224 39.433 ;
 RECT 14.336 37.973 14.392 38.173 ;
 RECT 14.168 37.973 14.224 38.173 ;
 RECT 13.664 39.367 13.72 39.567 ;
 RECT 15.008 39.443 15.064 39.643 ;
 RECT 14.84 39.917 14.896 40.082 ;
 RECT 14.672 39.917 14.728 40.082 ;
 RECT 13.664 38.107 13.72 38.307 ;
 RECT 15.008 38.183 15.064 38.383 ;
 RECT 14.84 38.657 14.896 38.822 ;
 RECT 14.672 38.657 14.728 38.822 ;
 RECT 13.664 36.847 13.72 37.047 ;
 RECT 15.008 36.923 15.064 37.123 ;
 RECT 14.84 37.397 14.896 37.562 ;
 RECT 14.672 37.397 14.728 37.562 ;
 RECT 13.664 35.587 13.72 35.787 ;
 RECT 15.008 35.663 15.064 35.863 ;
 RECT 14.84 36.137 14.896 36.302 ;
 RECT 14.672 36.137 14.728 36.302 ;
 RECT 15.176 36.3635 15.232 36.5635 ;
 RECT 12.824 36.148 12.88 36.348 ;
 RECT 13.496 36.159 13.552 36.359 ;
 RECT 13.328 36.097 13.384 36.297 ;
 RECT 13.16 36.148 13.216 36.348 ;
 RECT 12.488 36.178 12.544 36.378 ;
 RECT 12.992 36.148 13.048 36.348 ;
 RECT 12.656 36.178 12.712 36.378 ;
 END
 END vss.gds2960
 PIN vss.gds2961
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 39.96 15.418 40.16 ;
 END
 END vss.gds2961
 PIN vss.gds2962
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.438 38.8595 17.494 39.0595 ;
 END
 END vss.gds2962
 PIN vss.gds2963
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 38.0475 20.274 38.2475 ;
 END
 END vss.gds2963
 PIN vss.gds2964
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.702 36.2835 18.762 36.4835 ;
 END
 END vss.gds2964
 PIN vss.gds2965
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 39.217 16.146 39.417 ;
 END
 END vss.gds2965
 PIN vss.gds2966
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.038 36.2835 19.098 36.4835 ;
 END
 END vss.gds2966
 PIN vss.gds2967
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.206 36.2835 19.266 36.4835 ;
 END
 END vss.gds2967
 PIN vss.gds2968
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.374 36.2835 19.434 36.4835 ;
 END
 END vss.gds2968
 PIN vss.gds2969
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 37.957 16.146 38.157 ;
 END
 END vss.gds2969
 PIN vss.gds2970
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.71 36.2835 19.77 36.4835 ;
 END
 END vss.gds2970
 PIN vss.gds2971
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 36.697 16.146 36.897 ;
 END
 END vss.gds2971
 PIN vss.gds2972
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.878 36.2835 19.938 36.4835 ;
 END
 END vss.gds2972
 PIN vss.gds2973
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.534 36.2835 18.594 36.4835 ;
 END
 END vss.gds2973
 PIN vss.gds2974
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 36.756 16.814 36.956 ;
 END
 END vss.gds2974
 PIN vss.gds2975
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.366 36.2835 18.426 36.4835 ;
 END
 END vss.gds2975
 PIN vss.gds2976
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 39.839 17.314 40.039 ;
 END
 END vss.gds2976
 PIN vss.gds2977
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.986 36.067 18.026 36.267 ;
 END
 END vss.gds2977
 PIN vss.gds2978
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 38.0475 18.93 38.2475 ;
 END
 END vss.gds2978
 PIN vss.gds2979
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 38.0475 19.602 38.2475 ;
 END
 END vss.gds2979
 PIN vss.gds2980
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 38.0065 16.994 38.2065 ;
 END
 END vss.gds2980
 PIN vss.gds2981
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.046 36.2835 20.106 36.4835 ;
 END
 END vss.gds2981
 PIN vss.gds2982
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 38.088 15.842 38.288 ;
 END
 END vss.gds2982
 PIN vss.gds2983
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 37.885 18.258 38.085 ;
 END
 END vss.gds2983
 PIN vss.gds2984
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 38.2035 17.834 38.4035 ;
 END
 END vss.gds2984
 PIN vss.gds2985
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 38.1905 16.49 38.3905 ;
 END
 END vss.gds2985
 PIN vss.gds2986
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 16.52 36.14 16.576 36.293 ;
 RECT 15.764 36.137 15.82 36.302 ;
 RECT 15.596 36.137 15.652 36.302 ;
 RECT 15.596 36.364 15.652 36.564 ;
 RECT 15.848 36.367 15.904 36.567 ;
 RECT 16.52 37.4 16.576 37.553 ;
 RECT 15.764 37.397 15.82 37.562 ;
 RECT 15.596 37.397 15.652 37.562 ;
 RECT 15.596 37.624 15.652 37.824 ;
 RECT 15.848 37.627 15.904 37.827 ;
 RECT 16.52 38.66 16.576 38.813 ;
 RECT 15.764 38.657 15.82 38.822 ;
 RECT 15.596 38.657 15.652 38.822 ;
 RECT 15.596 38.884 15.652 39.084 ;
 RECT 15.848 38.887 15.904 39.087 ;
 RECT 16.52 39.92 16.576 40.073 ;
 RECT 15.764 39.917 15.82 40.082 ;
 RECT 15.596 39.917 15.652 40.082 ;
 RECT 15.596 40.144 15.652 40.344 ;
 RECT 15.848 40.147 15.904 40.347 ;
 RECT 16.352 39.5435 16.408 39.7435 ;
 RECT 16.856 39.2915 16.912 39.4915 ;
 RECT 16.856 38.0315 16.912 38.2315 ;
 RECT 16.352 38.2835 16.408 38.4835 ;
 RECT 16.352 37.0235 16.408 37.2235 ;
 RECT 16.856 36.7715 16.912 36.9715 ;
 RECT 16.352 35.7635 16.408 35.9635 ;
 RECT 16.856 35.5115 16.912 35.7115 ;
 RECT 15.428 39.443 15.484 39.643 ;
 RECT 15.428 38.183 15.484 38.383 ;
 RECT 15.428 36.923 15.484 37.123 ;
 RECT 15.428 35.663 15.484 35.863 ;
 RECT 17.864 36.178 17.92 36.378 ;
 RECT 17.696 36.1855 17.752 36.3855 ;
 RECT 17.528 36.178 17.584 36.378 ;
 RECT 17.36 36.178 17.416 36.378 ;
 RECT 17.192 36.178 17.248 36.378 ;
 RECT 18.032 36.178 18.088 36.378 ;
 RECT 17.024 36.293 17.08 36.493 ;
 END
 END vss.gds2986
 PIN vss.gds2987
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.17 36.2835 25.23 36.4835 ;
 END
 END vss.gds2987
 PIN vss.gds2988
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.002 36.2835 25.062 36.4835 ;
 END
 END vss.gds2988
 PIN vss.gds2989
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.834 36.2835 24.894 36.4835 ;
 END
 END vss.gds2989
 PIN vss.gds2990
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.498 36.2835 24.558 36.4835 ;
 END
 END vss.gds2990
 PIN vss.gds2991
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.33 36.2835 24.39 36.4835 ;
 END
 END vss.gds2991
 PIN vss.gds2992
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.162 36.2835 24.222 36.4835 ;
 END
 END vss.gds2992
 PIN vss.gds2993
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.382 36.2835 20.442 36.4835 ;
 END
 END vss.gds2993
 PIN vss.gds2994
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.55 36.2835 20.61 36.4835 ;
 END
 END vss.gds2994
 PIN vss.gds2995
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.718 36.2835 20.778 36.4835 ;
 END
 END vss.gds2995
 PIN vss.gds2996
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.054 36.2835 21.114 36.4835 ;
 END
 END vss.gds2996
 PIN vss.gds2997
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.222 36.2835 21.282 36.4835 ;
 END
 END vss.gds2997
 PIN vss.gds2998
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.39 36.2835 21.45 36.4835 ;
 END
 END vss.gds2998
 PIN vss.gds2999
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.726 36.2835 21.786 36.4835 ;
 END
 END vss.gds2999
 PIN vss.gds3000
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.894 36.2835 21.954 36.4835 ;
 END
 END vss.gds3000
 PIN vss.gds3001
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.062 36.2835 22.122 36.4835 ;
 END
 END vss.gds3001
 PIN vss.gds3002
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 38.0475 24.726 38.2475 ;
 END
 END vss.gds3002
 PIN vss.gds3003
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 38.0475 21.618 38.2475 ;
 END
 END vss.gds3003
 PIN vss.gds3004
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 38.0475 20.946 38.2475 ;
 END
 END vss.gds3004
 PIN vss.gds3005
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 38.0475 22.29 38.2475 ;
 END
 END vss.gds3005
 PIN vss.gds3006
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.398 36.2835 22.458 36.4835 ;
 END
 END vss.gds3006
 PIN vss.gds3007
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.566 36.2835 22.626 36.4835 ;
 END
 END vss.gds3007
 PIN vss.gds3008
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.734 36.2835 22.794 36.4835 ;
 END
 END vss.gds3008
 PIN vss.gds3009
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.07 36.2835 23.13 36.4835 ;
 END
 END vss.gds3009
 PIN vss.gds3010
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.238 36.2835 23.298 36.4835 ;
 END
 END vss.gds3010
 PIN vss.gds3011
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.406 36.2835 23.466 36.4835 ;
 END
 END vss.gds3011
 PIN vss.gds3012
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 38.0475 22.962 38.2475 ;
 END
 END vss.gds3012
 PIN vss.gds3013
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 38.0475 23.634 38.2475 ;
 END
 END vss.gds3013
 PIN vss.gds3014
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 23.912 39.38 23.968 39.58 ;
 RECT 23.912 38.12 23.968 38.32 ;
 RECT 23.912 36.86 23.968 37.06 ;
 RECT 23.912 35.6 23.968 35.8 ;
 RECT 23.744 38.05 23.8 38.25 ;
 END
 END vss.gds3014
 PIN vss.gds3015
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.202 36.2835 29.262 36.4835 ;
 END
 END vss.gds3015
 PIN vss.gds3016
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.034 36.2835 29.094 36.4835 ;
 END
 END vss.gds3016
 PIN vss.gds3017
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.866 36.2835 28.926 36.4835 ;
 END
 END vss.gds3017
 PIN vss.gds3018
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.53 36.2835 28.59 36.4835 ;
 END
 END vss.gds3018
 PIN vss.gds3019
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.362 36.2835 28.422 36.4835 ;
 END
 END vss.gds3019
 PIN vss.gds3020
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.194 36.2835 28.254 36.4835 ;
 END
 END vss.gds3020
 PIN vss.gds3021
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.858 36.2835 27.918 36.4835 ;
 END
 END vss.gds3021
 PIN vss.gds3022
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.69 36.2835 27.75 36.4835 ;
 END
 END vss.gds3022
 PIN vss.gds3023
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.522 36.2835 27.582 36.4835 ;
 END
 END vss.gds3023
 PIN vss.gds3024
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.186 36.2835 27.246 36.4835 ;
 END
 END vss.gds3024
 PIN vss.gds3025
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.018 36.2835 27.078 36.4835 ;
 END
 END vss.gds3025
 PIN vss.gds3026
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.85 36.2835 26.91 36.4835 ;
 END
 END vss.gds3026
 PIN vss.gds3027
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.514 36.2835 26.574 36.4835 ;
 END
 END vss.gds3027
 PIN vss.gds3028
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.346 36.2835 26.406 36.4835 ;
 END
 END vss.gds3028
 PIN vss.gds3029
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.178 36.2835 26.238 36.4835 ;
 END
 END vss.gds3029
 PIN vss.gds3030
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.842 36.2835 25.902 36.4835 ;
 END
 END vss.gds3030
 PIN vss.gds3031
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.674 36.2835 25.734 36.4835 ;
 END
 END vss.gds3031
 PIN vss.gds3032
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.506 36.2835 25.566 36.4835 ;
 END
 END vss.gds3032
 PIN vss.gds3033
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 38.0475 28.758 38.2475 ;
 END
 END vss.gds3033
 PIN vss.gds3034
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 38.0475 28.086 38.2475 ;
 END
 END vss.gds3034
 PIN vss.gds3035
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 38.0475 27.414 38.2475 ;
 END
 END vss.gds3035
 PIN vss.gds3036
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 38.0475 26.742 38.2475 ;
 END
 END vss.gds3036
 PIN vss.gds3037
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 38.0475 26.07 38.2475 ;
 END
 END vss.gds3037
 PIN vss.gds3038
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 38.0475 25.398 38.2475 ;
 END
 END vss.gds3038
 PIN vss.gds3039
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 37.885 29.43 38.085 ;
 END
 END vss.gds3039
 PIN vss.gds3040
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 36.9695 30.11 37.1695 ;
 END
 END vss.gds3040
 PIN vss.gds3041
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 38.2035 29.87 38.4035 ;
 END
 END vss.gds3041
 PIN vss.gds3042
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 38.587 29.642 38.787 ;
 END
 END vss.gds3042
 PIN vss.gds3043
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.876 36.148 29.932 36.348 ;
 RECT 29.708 36.178 29.764 36.378 ;
 RECT 30.212 36.148 30.268 36.348 ;
 RECT 29.54 36.178 29.596 36.378 ;
 RECT 30.044 36.148 30.1 36.348 ;
 END
 END vss.gds3043
 PIN vss.gds3044
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 37.242 31.922 37.442 ;
 END
 END vss.gds3044
 PIN vss.gds3045
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 37.202 30.95 37.402 ;
 END
 END vss.gds3045
 PIN vss.gds3046
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 35.942 30.95 36.142 ;
 END
 END vss.gds3046
 PIN vss.gds3047
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 35.982 31.922 36.182 ;
 END
 END vss.gds3047
 PIN vss.gds3048
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 39.762 31.922 39.962 ;
 END
 END vss.gds3048
 PIN vss.gds3049
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 38.502 31.922 38.702 ;
 END
 END vss.gds3049
 PIN vss.gds3050
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 39.722 30.95 39.922 ;
 END
 END vss.gds3050
 PIN vss.gds3051
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.314 39.276 30.37 39.476 ;
 END
 END vss.gds3051
 PIN vss.gds3052
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.49 38.8595 34.546 39.0595 ;
 END
 END vss.gds3052
 PIN vss.gds3053
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 39.217 33.198 39.417 ;
 END
 END vss.gds3053
 PIN vss.gds3054
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 37.957 33.198 38.157 ;
 END
 END vss.gds3054
 PIN vss.gds3055
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 36.697 33.198 36.897 ;
 END
 END vss.gds3055
 PIN vss.gds3056
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 36.756 33.866 36.956 ;
 END
 END vss.gds3056
 PIN vss.gds3057
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 38.462 30.95 38.662 ;
 END
 END vss.gds3057
 PIN vss.gds3058
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 38.088 32.214 38.288 ;
 END
 END vss.gds3058
 PIN vss.gds3059
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 38.0065 34.046 38.2065 ;
 END
 END vss.gds3059
 PIN vss.gds3060
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 39.839 34.366 40.039 ;
 END
 END vss.gds3060
 PIN vss.gds3061
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 39.96 32.47 40.16 ;
 END
 END vss.gds3061
 PIN vss.gds3062
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.038 36.067 35.078 36.267 ;
 END
 END vss.gds3062
 PIN vss.gds3063
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 38.0475 30.71 38.2475 ;
 END
 END vss.gds3063
 PIN vss.gds3064
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 38.088 32.894 38.288 ;
 END
 END vss.gds3064
 PIN vss.gds3065
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 38.1905 33.542 38.3905 ;
 END
 END vss.gds3065
 PIN vss.gds3066
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 38.088 31.55 38.288 ;
 END
 END vss.gds3066
 PIN vss.gds3067
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 38.2035 34.886 38.4035 ;
 END
 END vss.gds3067
 PIN vss.gds3068
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 33.572 36.14 33.628 36.293 ;
 RECT 31.052 36.12 31.108 36.293 ;
 RECT 31.22 36.093 31.276 36.293 ;
 RECT 32.816 36.137 32.872 36.302 ;
 RECT 32.648 36.137 32.704 36.302 ;
 RECT 31.892 36.137 31.948 36.302 ;
 RECT 31.724 36.137 31.78 36.302 ;
 RECT 33.572 37.4 33.628 37.553 ;
 RECT 31.052 37.38 31.108 37.553 ;
 RECT 31.22 37.353 31.276 37.553 ;
 RECT 32.816 37.397 32.872 37.562 ;
 RECT 32.648 37.397 32.704 37.562 ;
 RECT 31.892 37.397 31.948 37.562 ;
 RECT 31.724 37.397 31.78 37.562 ;
 RECT 33.572 38.66 33.628 38.813 ;
 RECT 31.052 38.64 31.108 38.813 ;
 RECT 31.22 38.613 31.276 38.813 ;
 RECT 32.816 38.657 32.872 38.822 ;
 RECT 32.648 38.657 32.704 38.822 ;
 RECT 31.892 38.657 31.948 38.822 ;
 RECT 31.724 38.657 31.78 38.822 ;
 RECT 33.572 39.92 33.628 40.073 ;
 RECT 31.052 39.9 31.108 40.073 ;
 RECT 31.22 39.873 31.276 40.073 ;
 RECT 32.816 39.917 32.872 40.082 ;
 RECT 32.648 39.917 32.704 40.082 ;
 RECT 31.892 39.917 31.948 40.082 ;
 RECT 31.724 39.917 31.78 40.082 ;
 RECT 32.648 36.364 32.704 36.564 ;
 RECT 32.9 36.367 32.956 36.567 ;
 RECT 32.648 37.624 32.704 37.824 ;
 RECT 32.9 37.627 32.956 37.827 ;
 RECT 32.648 40.144 32.704 40.344 ;
 RECT 32.9 40.147 32.956 40.347 ;
 RECT 32.648 38.884 32.704 39.084 ;
 RECT 32.9 38.887 32.956 39.087 ;
 RECT 31.388 37.973 31.444 38.173 ;
 RECT 31.22 37.973 31.276 38.173 ;
 RECT 32.06 38.183 32.116 38.383 ;
 RECT 32.48 38.183 32.536 38.383 ;
 RECT 30.716 38.107 30.772 38.307 ;
 RECT 33.404 38.2835 33.46 38.4835 ;
 RECT 33.908 38.0315 33.964 38.2315 ;
 RECT 33.908 39.2915 33.964 39.4915 ;
 RECT 33.404 39.5435 33.46 39.7435 ;
 RECT 32.06 39.443 32.116 39.643 ;
 RECT 32.48 39.443 32.536 39.643 ;
 RECT 31.388 39.233 31.444 39.433 ;
 RECT 31.22 39.233 31.276 39.433 ;
 RECT 30.716 39.367 30.772 39.567 ;
 RECT 33.908 36.7715 33.964 36.9715 ;
 RECT 33.404 37.0235 33.46 37.2235 ;
 RECT 32.06 36.923 32.116 37.123 ;
 RECT 32.48 36.923 32.536 37.123 ;
 RECT 31.388 36.713 31.444 36.913 ;
 RECT 31.22 36.713 31.276 36.913 ;
 RECT 30.716 36.847 30.772 37.047 ;
 RECT 33.908 35.5115 33.964 35.7115 ;
 RECT 33.404 35.7635 33.46 35.9635 ;
 RECT 32.06 35.663 32.116 35.863 ;
 RECT 32.48 35.663 32.536 35.863 ;
 RECT 31.388 35.453 31.444 35.653 ;
 RECT 31.22 35.453 31.276 35.653 ;
 RECT 30.716 35.587 30.772 35.787 ;
 RECT 30.548 36.159 30.604 36.359 ;
 RECT 34.916 36.178 34.972 36.378 ;
 RECT 32.228 36.3635 32.284 36.5635 ;
 RECT 30.38 36.097 30.436 36.297 ;
 RECT 34.748 36.1855 34.804 36.3855 ;
 RECT 34.58 36.178 34.636 36.378 ;
 RECT 34.412 36.178 34.468 36.378 ;
 RECT 34.244 36.178 34.3 36.378 ;
 RECT 34.076 36.293 34.132 36.493 ;
 RECT 35.084 36.178 35.14 36.378 ;
 END
 END vss.gds3068
 PIN vss.gds3069
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.122 36.2835 40.182 36.4835 ;
 END
 END vss.gds3069
 PIN vss.gds3070
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.754 36.2835 35.814 36.4835 ;
 END
 END vss.gds3070
 PIN vss.gds3071
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.09 36.2835 36.15 36.4835 ;
 END
 END vss.gds3071
 PIN vss.gds3072
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.258 36.2835 36.318 36.4835 ;
 END
 END vss.gds3072
 PIN vss.gds3073
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.426 36.2835 36.486 36.4835 ;
 END
 END vss.gds3073
 PIN vss.gds3074
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 38.0475 36.654 38.2475 ;
 END
 END vss.gds3074
 PIN vss.gds3075
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.762 36.2835 36.822 36.4835 ;
 END
 END vss.gds3075
 PIN vss.gds3076
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.93 36.2835 36.99 36.4835 ;
 END
 END vss.gds3076
 PIN vss.gds3077
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.098 36.2835 37.158 36.4835 ;
 END
 END vss.gds3077
 PIN vss.gds3078
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 38.0475 37.326 38.2475 ;
 END
 END vss.gds3078
 PIN vss.gds3079
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.434 36.2835 37.494 36.4835 ;
 END
 END vss.gds3079
 PIN vss.gds3080
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.602 36.2835 37.662 36.4835 ;
 END
 END vss.gds3080
 PIN vss.gds3081
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.77 36.2835 37.83 36.4835 ;
 END
 END vss.gds3081
 PIN vss.gds3082
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 38.0475 37.998 38.2475 ;
 END
 END vss.gds3082
 PIN vss.gds3083
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.106 36.2835 38.166 36.4835 ;
 END
 END vss.gds3083
 PIN vss.gds3084
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.274 36.2835 38.334 36.4835 ;
 END
 END vss.gds3084
 PIN vss.gds3085
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.442 36.2835 38.502 36.4835 ;
 END
 END vss.gds3085
 PIN vss.gds3086
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.778 36.2835 38.838 36.4835 ;
 END
 END vss.gds3086
 PIN vss.gds3087
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.946 36.2835 39.006 36.4835 ;
 END
 END vss.gds3087
 PIN vss.gds3088
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.45 36.2835 39.51 36.4835 ;
 END
 END vss.gds3088
 PIN vss.gds3089
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.618 36.2835 39.678 36.4835 ;
 END
 END vss.gds3089
 PIN vss.gds3090
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.586 36.2835 35.646 36.4835 ;
 END
 END vss.gds3090
 PIN vss.gds3091
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.786 36.2835 39.846 36.4835 ;
 END
 END vss.gds3091
 PIN vss.gds3092
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.114 36.2835 39.174 36.4835 ;
 END
 END vss.gds3092
 PIN vss.gds3093
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.418 36.2835 35.478 36.4835 ;
 END
 END vss.gds3093
 PIN vss.gds3094
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 38.0475 38.67 38.2475 ;
 END
 END vss.gds3094
 PIN vss.gds3095
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 38.0475 35.982 38.2475 ;
 END
 END vss.gds3095
 PIN vss.gds3096
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 38.0475 40.014 38.2475 ;
 END
 END vss.gds3096
 PIN vss.gds3097
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 37.885 35.31 38.085 ;
 END
 END vss.gds3097
 PIN vss.gds3098
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 38.0475 39.342 38.2475 ;
 END
 END vss.gds3098
 PIN vss.gds3099
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 38.0475 45.138 38.2475 ;
 END
 END vss.gds3099
 PIN vss.gds3100
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.91 36.2835 44.97 36.4835 ;
 END
 END vss.gds3100
 PIN vss.gds3101
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.742 36.2835 44.802 36.4835 ;
 END
 END vss.gds3101
 PIN vss.gds3102
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.574 36.2835 44.634 36.4835 ;
 END
 END vss.gds3102
 PIN vss.gds3103
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 38.0475 44.466 38.2475 ;
 END
 END vss.gds3103
 PIN vss.gds3104
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.238 36.2835 44.298 36.4835 ;
 END
 END vss.gds3104
 PIN vss.gds3105
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.07 36.2835 44.13 36.4835 ;
 END
 END vss.gds3105
 PIN vss.gds3106
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.902 36.2835 43.962 36.4835 ;
 END
 END vss.gds3106
 PIN vss.gds3107
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 38.0475 43.794 38.2475 ;
 END
 END vss.gds3107
 PIN vss.gds3108
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.566 36.2835 43.626 36.4835 ;
 END
 END vss.gds3108
 PIN vss.gds3109
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.398 36.2835 43.458 36.4835 ;
 END
 END vss.gds3109
 PIN vss.gds3110
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.23 36.2835 43.29 36.4835 ;
 END
 END vss.gds3110
 PIN vss.gds3111
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 38.0475 43.122 38.2475 ;
 END
 END vss.gds3111
 PIN vss.gds3112
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.894 36.2835 42.954 36.4835 ;
 END
 END vss.gds3112
 PIN vss.gds3113
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.726 36.2835 42.786 36.4835 ;
 END
 END vss.gds3113
 PIN vss.gds3114
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.558 36.2835 42.618 36.4835 ;
 END
 END vss.gds3114
 PIN vss.gds3115
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 38.0475 42.45 38.2475 ;
 END
 END vss.gds3115
 PIN vss.gds3116
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.222 36.2835 42.282 36.4835 ;
 END
 END vss.gds3116
 PIN vss.gds3117
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.054 36.2835 42.114 36.4835 ;
 END
 END vss.gds3117
 PIN vss.gds3118
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.886 36.2835 41.946 36.4835 ;
 END
 END vss.gds3118
 PIN vss.gds3119
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 38.0475 41.778 38.2475 ;
 END
 END vss.gds3119
 PIN vss.gds3120
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.55 36.2835 41.61 36.4835 ;
 END
 END vss.gds3120
 PIN vss.gds3121
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.382 36.2835 41.442 36.4835 ;
 END
 END vss.gds3121
 PIN vss.gds3122
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.214 36.2835 41.274 36.4835 ;
 END
 END vss.gds3122
 PIN vss.gds3123
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.29 36.2835 40.35 36.4835 ;
 END
 END vss.gds3123
 PIN vss.gds3124
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.458 36.2835 40.518 36.4835 ;
 END
 END vss.gds3124
 PIN vss.gds3125
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 38.0475 40.686 38.2475 ;
 END
 END vss.gds3125
 PIN vss.gds3126
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 40.964 38.12 41.02 38.32 ;
 RECT 40.964 39.38 41.02 39.58 ;
 RECT 40.964 36.86 41.02 37.06 ;
 RECT 40.964 35.6 41.02 35.8 ;
 RECT 40.796 38.05 40.852 38.25 ;
 END
 END vss.gds3126
 PIN vss.gds3127
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 37.242 48.974 37.442 ;
 END
 END vss.gds3127
 PIN vss.gds3128
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 35.982 48.974 36.182 ;
 END
 END vss.gds3128
 PIN vss.gds3129
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 39.762 48.974 39.962 ;
 END
 END vss.gds3129
 PIN vss.gds3130
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 38.502 48.974 38.702 ;
 END
 END vss.gds3130
 PIN vss.gds3131
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 35.942 48.002 36.142 ;
 END
 END vss.gds3131
 PIN vss.gds3132
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 37.202 48.002 37.402 ;
 END
 END vss.gds3132
 PIN vss.gds3133
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 39.722 48.002 39.922 ;
 END
 END vss.gds3133
 PIN vss.gds3134
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.366 39.276 47.422 39.476 ;
 END
 END vss.gds3134
 PIN vss.gds3135
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 37.885 46.482 38.085 ;
 END
 END vss.gds3135
 PIN vss.gds3136
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.254 36.2835 46.314 36.4835 ;
 END
 END vss.gds3136
 PIN vss.gds3137
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.086 36.2835 46.146 36.4835 ;
 END
 END vss.gds3137
 PIN vss.gds3138
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.918 36.2835 45.978 36.4835 ;
 END
 END vss.gds3138
 PIN vss.gds3139
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 38.0475 45.81 38.2475 ;
 END
 END vss.gds3139
 PIN vss.gds3140
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.582 36.2835 45.642 36.4835 ;
 END
 END vss.gds3140
 PIN vss.gds3141
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.414 36.2835 45.474 36.4835 ;
 END
 END vss.gds3141
 PIN vss.gds3142
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.246 36.2835 45.306 36.4835 ;
 END
 END vss.gds3142
 PIN vss.gds3143
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 36.9695 47.162 37.1695 ;
 END
 END vss.gds3143
 PIN vss.gds3144
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 39.96 49.522 40.16 ;
 END
 END vss.gds3144
 PIN vss.gds3145
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 39.217 50.25 39.417 ;
 END
 END vss.gds3145
 PIN vss.gds3146
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 37.957 50.25 38.157 ;
 END
 END vss.gds3146
 PIN vss.gds3147
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 36.697 50.25 36.897 ;
 END
 END vss.gds3147
 PIN vss.gds3148
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 38.462 48.002 38.662 ;
 END
 END vss.gds3148
 PIN vss.gds3149
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 38.2035 46.922 38.4035 ;
 END
 END vss.gds3149
 PIN vss.gds3150
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 38.587 46.694 38.787 ;
 END
 END vss.gds3150
 PIN vss.gds3151
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 38.0475 47.762 38.2475 ;
 END
 END vss.gds3151
 PIN vss.gds3152
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 38.088 49.266 38.288 ;
 END
 END vss.gds3152
 PIN vss.gds3153
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 38.088 48.602 38.288 ;
 END
 END vss.gds3153
 PIN vss.gds3154
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 38.088 49.946 38.288 ;
 END
 END vss.gds3154
 PIN vss.gds3155
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 48.104 36.12 48.16 36.293 ;
 RECT 48.272 36.093 48.328 36.293 ;
 RECT 49.868 36.137 49.924 36.302 ;
 RECT 49.7 36.137 49.756 36.302 ;
 RECT 48.944 36.137 49 36.302 ;
 RECT 48.776 36.137 48.832 36.302 ;
 RECT 48.104 37.38 48.16 37.553 ;
 RECT 48.272 37.353 48.328 37.553 ;
 RECT 49.868 37.397 49.924 37.562 ;
 RECT 49.7 37.397 49.756 37.562 ;
 RECT 48.944 37.397 49 37.562 ;
 RECT 48.776 37.397 48.832 37.562 ;
 RECT 48.104 38.64 48.16 38.813 ;
 RECT 48.272 38.613 48.328 38.813 ;
 RECT 49.868 38.657 49.924 38.822 ;
 RECT 49.7 38.657 49.756 38.822 ;
 RECT 48.944 38.657 49 38.822 ;
 RECT 48.776 38.657 48.832 38.822 ;
 RECT 48.104 39.9 48.16 40.073 ;
 RECT 48.272 39.873 48.328 40.073 ;
 RECT 49.868 39.917 49.924 40.082 ;
 RECT 49.7 39.917 49.756 40.082 ;
 RECT 48.944 39.917 49 40.082 ;
 RECT 48.776 39.917 48.832 40.082 ;
 RECT 49.7 36.364 49.756 36.564 ;
 RECT 49.952 36.367 50.008 36.567 ;
 RECT 49.7 38.884 49.756 39.084 ;
 RECT 49.952 38.887 50.008 39.087 ;
 RECT 49.7 40.144 49.756 40.344 ;
 RECT 49.952 40.147 50.008 40.347 ;
 RECT 49.7 37.624 49.756 37.824 ;
 RECT 49.952 37.627 50.008 37.827 ;
 RECT 48.44 37.973 48.496 38.173 ;
 RECT 48.272 37.973 48.328 38.173 ;
 RECT 49.112 38.183 49.168 38.383 ;
 RECT 49.532 38.183 49.588 38.383 ;
 RECT 49.112 39.443 49.168 39.643 ;
 RECT 49.532 39.443 49.588 39.643 ;
 RECT 48.44 39.233 48.496 39.433 ;
 RECT 48.272 39.233 48.328 39.433 ;
 RECT 47.768 39.367 47.824 39.567 ;
 RECT 47.768 38.107 47.824 38.307 ;
 RECT 49.112 36.923 49.168 37.123 ;
 RECT 49.532 36.923 49.588 37.123 ;
 RECT 48.44 36.713 48.496 36.913 ;
 RECT 48.272 36.713 48.328 36.913 ;
 RECT 47.768 36.847 47.824 37.047 ;
 RECT 49.112 35.663 49.168 35.863 ;
 RECT 49.532 35.663 49.588 35.863 ;
 RECT 48.44 35.453 48.496 35.653 ;
 RECT 48.272 35.453 48.328 35.653 ;
 RECT 47.768 35.587 47.824 35.787 ;
 RECT 47.6 36.159 47.656 36.359 ;
 RECT 49.28 36.3635 49.336 36.5635 ;
 RECT 46.928 36.148 46.984 36.348 ;
 RECT 47.432 36.097 47.488 36.297 ;
 RECT 47.264 36.148 47.32 36.348 ;
 RECT 46.592 36.178 46.648 36.378 ;
 RECT 46.76 36.178 46.816 36.378 ;
 RECT 47.096 36.148 47.152 36.348 ;
 END
 END vss.gds3155
 PIN vss.gds3156
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.542 38.8595 51.598 39.0595 ;
 END
 END vss.gds3156
 PIN vss.gds3157
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 36.756 50.918 36.956 ;
 END
 END vss.gds3157
 PIN vss.gds3158
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.638 36.2835 52.698 36.4835 ;
 END
 END vss.gds3158
 PIN vss.gds3159
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.806 36.2835 52.866 36.4835 ;
 END
 END vss.gds3159
 PIN vss.gds3160
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.142 36.2835 53.202 36.4835 ;
 END
 END vss.gds3160
 PIN vss.gds3161
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.31 36.2835 53.37 36.4835 ;
 END
 END vss.gds3161
 PIN vss.gds3162
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.478 36.2835 53.538 36.4835 ;
 END
 END vss.gds3162
 PIN vss.gds3163
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.814 36.2835 53.874 36.4835 ;
 END
 END vss.gds3163
 PIN vss.gds3164
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.982 36.2835 54.042 36.4835 ;
 END
 END vss.gds3164
 PIN vss.gds3165
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.15 36.2835 54.21 36.4835 ;
 END
 END vss.gds3165
 PIN vss.gds3166
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.486 36.2835 54.546 36.4835 ;
 END
 END vss.gds3166
 PIN vss.gds3167
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.654 36.2835 54.714 36.4835 ;
 END
 END vss.gds3167
 PIN vss.gds3168
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.822 36.2835 54.882 36.4835 ;
 END
 END vss.gds3168
 PIN vss.gds3169
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 38.0475 55.05 38.2475 ;
 END
 END vss.gds3169
 PIN vss.gds3170
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.158 36.2835 55.218 36.4835 ;
 END
 END vss.gds3170
 PIN vss.gds3171
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 38.0475 54.378 38.2475 ;
 END
 END vss.gds3171
 PIN vss.gds3172
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 38.0475 53.706 38.2475 ;
 END
 END vss.gds3172
 PIN vss.gds3173
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.47 36.2835 52.53 36.4835 ;
 END
 END vss.gds3173
 PIN vss.gds3174
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 39.839 51.418 40.039 ;
 END
 END vss.gds3174
 PIN vss.gds3175
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.09 36.067 52.13 36.267 ;
 END
 END vss.gds3175
 PIN vss.gds3176
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 38.0065 51.098 38.2065 ;
 END
 END vss.gds3176
 PIN vss.gds3177
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 38.0475 53.034 38.2475 ;
 END
 END vss.gds3177
 PIN vss.gds3178
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 38.2035 51.938 38.4035 ;
 END
 END vss.gds3178
 PIN vss.gds3179
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 38.1905 50.594 38.3905 ;
 END
 END vss.gds3179
 PIN vss.gds3180
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 37.885 52.362 38.085 ;
 END
 END vss.gds3180
 PIN vss.gds3181
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 50.624 36.14 50.68 36.293 ;
 RECT 50.624 37.4 50.68 37.553 ;
 RECT 50.624 38.66 50.68 38.813 ;
 RECT 50.624 39.92 50.68 40.073 ;
 RECT 50.96 39.2915 51.016 39.4915 ;
 RECT 50.456 39.5435 50.512 39.7435 ;
 RECT 50.456 38.2835 50.512 38.4835 ;
 RECT 50.96 38.0315 51.016 38.2315 ;
 RECT 50.96 36.7715 51.016 36.9715 ;
 RECT 50.456 37.0235 50.512 37.2235 ;
 RECT 50.96 35.5115 51.016 35.7115 ;
 RECT 50.456 35.7635 50.512 35.9635 ;
 RECT 51.968 36.178 52.024 36.378 ;
 RECT 51.8 36.1855 51.856 36.3855 ;
 RECT 51.632 36.178 51.688 36.378 ;
 RECT 51.464 36.178 51.52 36.378 ;
 RECT 51.296 36.178 51.352 36.378 ;
 RECT 51.128 36.293 51.184 36.493 ;
 RECT 52.136 36.178 52.192 36.378 ;
 END
 END vss.gds3181
 PIN vss.gds3182
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 38.0475 60.174 38.2475 ;
 END
 END vss.gds3182
 PIN vss.gds3183
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.946 36.2835 60.006 36.4835 ;
 END
 END vss.gds3183
 PIN vss.gds3184
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.778 36.2835 59.838 36.4835 ;
 END
 END vss.gds3184
 PIN vss.gds3185
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.61 36.2835 59.67 36.4835 ;
 END
 END vss.gds3185
 PIN vss.gds3186
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 38.0475 59.502 38.2475 ;
 END
 END vss.gds3186
 PIN vss.gds3187
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.274 36.2835 59.334 36.4835 ;
 END
 END vss.gds3187
 PIN vss.gds3188
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.106 36.2835 59.166 36.4835 ;
 END
 END vss.gds3188
 PIN vss.gds3189
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.938 36.2835 58.998 36.4835 ;
 END
 END vss.gds3189
 PIN vss.gds3190
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 38.0475 58.83 38.2475 ;
 END
 END vss.gds3190
 PIN vss.gds3191
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.602 36.2835 58.662 36.4835 ;
 END
 END vss.gds3191
 PIN vss.gds3192
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.434 36.2835 58.494 36.4835 ;
 END
 END vss.gds3192
 PIN vss.gds3193
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.266 36.2835 58.326 36.4835 ;
 END
 END vss.gds3193
 PIN vss.gds3194
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.326 36.2835 55.386 36.4835 ;
 END
 END vss.gds3194
 PIN vss.gds3195
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.494 36.2835 55.554 36.4835 ;
 END
 END vss.gds3195
 PIN vss.gds3196
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.83 36.2835 55.89 36.4835 ;
 END
 END vss.gds3196
 PIN vss.gds3197
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.998 36.2835 56.058 36.4835 ;
 END
 END vss.gds3197
 PIN vss.gds3198
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.166 36.2835 56.226 36.4835 ;
 END
 END vss.gds3198
 PIN vss.gds3199
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.502 36.2835 56.562 36.4835 ;
 END
 END vss.gds3199
 PIN vss.gds3200
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.67 36.2835 56.73 36.4835 ;
 END
 END vss.gds3200
 PIN vss.gds3201
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.838 36.2835 56.898 36.4835 ;
 END
 END vss.gds3201
 PIN vss.gds3202
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.342 36.2835 57.402 36.4835 ;
 END
 END vss.gds3202
 PIN vss.gds3203
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.51 36.2835 57.57 36.4835 ;
 END
 END vss.gds3203
 PIN vss.gds3204
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 38.0475 55.722 38.2475 ;
 END
 END vss.gds3204
 PIN vss.gds3205
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 38.0475 56.394 38.2475 ;
 END
 END vss.gds3205
 PIN vss.gds3206
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.174 36.2835 57.234 36.4835 ;
 END
 END vss.gds3206
 PIN vss.gds3207
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 38.0475 57.738 38.2475 ;
 END
 END vss.gds3207
 PIN vss.gds3208
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 38.0475 57.066 38.2475 ;
 END
 END vss.gds3208
 PIN vss.gds3209
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 58.016 38.12 58.072 38.32 ;
 RECT 58.016 39.38 58.072 39.58 ;
 RECT 58.016 36.86 58.072 37.06 ;
 RECT 58.016 35.6 58.072 35.8 ;
 RECT 57.848 38.05 57.904 38.25 ;
 END
 END vss.gds3209
 PIN vss.gds3210
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 37.202 65.054 37.402 ;
 END
 END vss.gds3210
 PIN vss.gds3211
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 35.942 65.054 36.142 ;
 END
 END vss.gds3211
 PIN vss.gds3212
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 38.462 65.054 38.662 ;
 END
 END vss.gds3212
 PIN vss.gds3213
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 36.9695 64.214 37.1695 ;
 END
 END vss.gds3213
 PIN vss.gds3214
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.418 39.276 64.474 39.476 ;
 END
 END vss.gds3214
 PIN vss.gds3215
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 37.885 63.534 38.085 ;
 END
 END vss.gds3215
 PIN vss.gds3216
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.306 36.2835 63.366 36.4835 ;
 END
 END vss.gds3216
 PIN vss.gds3217
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.138 36.2835 63.198 36.4835 ;
 END
 END vss.gds3217
 PIN vss.gds3218
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.97 36.2835 63.03 36.4835 ;
 END
 END vss.gds3218
 PIN vss.gds3219
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 38.0475 62.862 38.2475 ;
 END
 END vss.gds3219
 PIN vss.gds3220
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.634 36.2835 62.694 36.4835 ;
 END
 END vss.gds3220
 PIN vss.gds3221
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.466 36.2835 62.526 36.4835 ;
 END
 END vss.gds3221
 PIN vss.gds3222
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.298 36.2835 62.358 36.4835 ;
 END
 END vss.gds3222
 PIN vss.gds3223
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 38.0475 62.19 38.2475 ;
 END
 END vss.gds3223
 PIN vss.gds3224
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.962 36.2835 62.022 36.4835 ;
 END
 END vss.gds3224
 PIN vss.gds3225
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.794 36.2835 61.854 36.4835 ;
 END
 END vss.gds3225
 PIN vss.gds3226
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.626 36.2835 61.686 36.4835 ;
 END
 END vss.gds3226
 PIN vss.gds3227
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 38.0475 61.518 38.2475 ;
 END
 END vss.gds3227
 PIN vss.gds3228
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.29 36.2835 61.35 36.4835 ;
 END
 END vss.gds3228
 PIN vss.gds3229
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.122 36.2835 61.182 36.4835 ;
 END
 END vss.gds3229
 PIN vss.gds3230
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.954 36.2835 61.014 36.4835 ;
 END
 END vss.gds3230
 PIN vss.gds3231
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 38.0475 60.846 38.2475 ;
 END
 END vss.gds3231
 PIN vss.gds3232
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.618 36.2835 60.678 36.4835 ;
 END
 END vss.gds3232
 PIN vss.gds3233
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.45 36.2835 60.51 36.4835 ;
 END
 END vss.gds3233
 PIN vss.gds3234
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.282 36.2835 60.342 36.4835 ;
 END
 END vss.gds3234
 PIN vss.gds3235
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 38.2035 63.974 38.4035 ;
 END
 END vss.gds3235
 PIN vss.gds3236
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 38.587 63.746 38.787 ;
 END
 END vss.gds3236
 PIN vss.gds3237
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 39.722 65.054 39.922 ;
 END
 END vss.gds3237
 PIN vss.gds3238
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 38.0475 64.814 38.2475 ;
 END
 END vss.gds3238
 PIN vss.gds3239
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 65.156 36.12 65.212 36.293 ;
 RECT 65.156 37.38 65.212 37.553 ;
 RECT 65.156 38.64 65.212 38.813 ;
 RECT 65.156 39.9 65.212 40.073 ;
 RECT 64.82 39.367 64.876 39.567 ;
 RECT 64.82 38.107 64.876 38.307 ;
 RECT 64.82 35.587 64.876 35.787 ;
 RECT 64.82 36.847 64.876 37.047 ;
 RECT 64.652 36.159 64.708 36.359 ;
 RECT 63.98 36.148 64.036 36.348 ;
 RECT 63.812 36.178 63.868 36.378 ;
 RECT 64.484 36.097 64.54 36.297 ;
 RECT 64.316 36.148 64.372 36.348 ;
 RECT 63.644 36.178 63.7 36.378 ;
 RECT 64.148 36.148 64.204 36.348 ;
 END
 END vss.gds3239
 PIN vss.gds3240
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 37.242 66.026 37.442 ;
 END
 END vss.gds3240
 PIN vss.gds3241
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 35.982 66.026 36.182 ;
 END
 END vss.gds3241
 PIN vss.gds3242
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 39.762 66.026 39.962 ;
 END
 END vss.gds3242
 PIN vss.gds3243
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 38.502 66.026 38.702 ;
 END
 END vss.gds3243
 PIN vss.gds3244
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 39.217 67.302 39.417 ;
 END
 END vss.gds3244
 PIN vss.gds3245
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 39.96 66.574 40.16 ;
 END
 END vss.gds3245
 PIN vss.gds3246
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.594 38.8595 68.65 39.0595 ;
 END
 END vss.gds3246
 PIN vss.gds3247
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 38.0065 68.15 38.2065 ;
 END
 END vss.gds3247
 PIN vss.gds3248
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.858 36.2835 69.918 36.4835 ;
 END
 END vss.gds3248
 PIN vss.gds3249
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.194 36.2835 70.254 36.4835 ;
 END
 END vss.gds3249
 PIN vss.gds3250
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.142 36.067 69.182 36.267 ;
 END
 END vss.gds3250
 PIN vss.gds3251
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 37.957 67.302 38.157 ;
 END
 END vss.gds3251
 PIN vss.gds3252
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 36.756 67.97 36.956 ;
 END
 END vss.gds3252
 PIN vss.gds3253
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 36.697 67.302 36.897 ;
 END
 END vss.gds3253
 PIN vss.gds3254
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.69 36.2835 69.75 36.4835 ;
 END
 END vss.gds3254
 PIN vss.gds3255
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 38.088 66.318 38.288 ;
 END
 END vss.gds3255
 PIN vss.gds3256
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.522 36.2835 69.582 36.4835 ;
 END
 END vss.gds3256
 PIN vss.gds3257
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 39.839 68.47 40.039 ;
 END
 END vss.gds3257
 PIN vss.gds3258
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 38.0475 70.086 38.2475 ;
 END
 END vss.gds3258
 PIN vss.gds3259
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 38.088 66.998 38.288 ;
 END
 END vss.gds3259
 PIN vss.gds3260
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 38.088 65.654 38.288 ;
 END
 END vss.gds3260
 PIN vss.gds3261
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 38.1905 67.646 38.3905 ;
 END
 END vss.gds3261
 PIN vss.gds3262
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 38.2035 68.99 38.4035 ;
 END
 END vss.gds3262
 PIN vss.gds3263
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 37.885 69.414 38.085 ;
 END
 END vss.gds3263
 PIN vss.gds3264
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 67.676 36.14 67.732 36.293 ;
 RECT 65.324 36.093 65.38 36.293 ;
 RECT 66.92 36.137 66.976 36.302 ;
 RECT 66.752 36.137 66.808 36.302 ;
 RECT 65.996 36.137 66.052 36.302 ;
 RECT 65.828 36.137 65.884 36.302 ;
 RECT 67.676 37.4 67.732 37.553 ;
 RECT 65.324 37.353 65.38 37.553 ;
 RECT 66.92 37.397 66.976 37.562 ;
 RECT 66.752 37.397 66.808 37.562 ;
 RECT 65.996 37.397 66.052 37.562 ;
 RECT 65.828 37.397 65.884 37.562 ;
 RECT 67.676 38.66 67.732 38.813 ;
 RECT 65.324 38.613 65.38 38.813 ;
 RECT 66.92 38.657 66.976 38.822 ;
 RECT 66.752 38.657 66.808 38.822 ;
 RECT 65.996 38.657 66.052 38.822 ;
 RECT 65.828 38.657 65.884 38.822 ;
 RECT 67.676 39.92 67.732 40.073 ;
 RECT 65.324 39.873 65.38 40.073 ;
 RECT 66.92 39.917 66.976 40.082 ;
 RECT 66.752 39.917 66.808 40.082 ;
 RECT 65.996 39.917 66.052 40.082 ;
 RECT 65.828 39.917 65.884 40.082 ;
 RECT 66.752 36.364 66.808 36.564 ;
 RECT 67.004 36.367 67.06 36.567 ;
 RECT 66.752 37.624 66.808 37.824 ;
 RECT 67.004 37.627 67.06 37.827 ;
 RECT 66.752 38.884 66.808 39.084 ;
 RECT 67.004 38.887 67.06 39.087 ;
 RECT 66.752 40.144 66.808 40.344 ;
 RECT 67.004 40.147 67.06 40.347 ;
 RECT 65.492 39.233 65.548 39.433 ;
 RECT 65.324 39.233 65.38 39.433 ;
 RECT 66.164 39.443 66.22 39.643 ;
 RECT 66.584 39.443 66.64 39.643 ;
 RECT 68.012 39.2915 68.068 39.4915 ;
 RECT 67.508 39.5435 67.564 39.7435 ;
 RECT 68.012 38.0315 68.068 38.2315 ;
 RECT 67.508 38.2835 67.564 38.4835 ;
 RECT 66.164 38.183 66.22 38.383 ;
 RECT 65.492 37.973 65.548 38.173 ;
 RECT 65.324 37.973 65.38 38.173 ;
 RECT 66.584 38.183 66.64 38.383 ;
 RECT 68.012 35.5115 68.068 35.7115 ;
 RECT 67.508 35.7635 67.564 35.9635 ;
 RECT 66.164 35.663 66.22 35.863 ;
 RECT 66.584 35.663 66.64 35.863 ;
 RECT 65.492 35.453 65.548 35.653 ;
 RECT 65.324 35.453 65.38 35.653 ;
 RECT 68.012 36.7715 68.068 36.9715 ;
 RECT 67.508 37.0235 67.564 37.2235 ;
 RECT 66.164 36.923 66.22 37.123 ;
 RECT 66.584 36.923 66.64 37.123 ;
 RECT 65.492 36.713 65.548 36.913 ;
 RECT 65.324 36.713 65.38 36.913 ;
 RECT 66.332 36.3635 66.388 36.5635 ;
 RECT 69.02 36.178 69.076 36.378 ;
 RECT 68.852 36.1855 68.908 36.3855 ;
 RECT 68.684 36.178 68.74 36.378 ;
 RECT 68.516 36.178 68.572 36.378 ;
 RECT 68.348 36.178 68.404 36.378 ;
 RECT 69.188 36.178 69.244 36.378 ;
 RECT 68.18 36.293 68.236 36.493 ;
 END
 END vss.gds3264
 PIN vss.gds3265
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.362 36.2835 70.422 36.4835 ;
 END
 END vss.gds3265
 PIN vss.gds3266
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.53 36.2835 70.59 36.4835 ;
 END
 END vss.gds3266
 PIN vss.gds3267
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.866 36.2835 70.926 36.4835 ;
 END
 END vss.gds3267
 PIN vss.gds3268
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.034 36.2835 71.094 36.4835 ;
 END
 END vss.gds3268
 PIN vss.gds3269
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.202 36.2835 71.262 36.4835 ;
 END
 END vss.gds3269
 PIN vss.gds3270
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 38.0475 71.43 38.2475 ;
 END
 END vss.gds3270
 PIN vss.gds3271
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.538 36.2835 71.598 36.4835 ;
 END
 END vss.gds3271
 PIN vss.gds3272
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.706 36.2835 71.766 36.4835 ;
 END
 END vss.gds3272
 PIN vss.gds3273
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.874 36.2835 71.934 36.4835 ;
 END
 END vss.gds3273
 PIN vss.gds3274
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 38.0475 72.102 38.2475 ;
 END
 END vss.gds3274
 PIN vss.gds3275
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.21 36.2835 72.27 36.4835 ;
 END
 END vss.gds3275
 PIN vss.gds3276
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.378 36.2835 72.438 36.4835 ;
 END
 END vss.gds3276
 PIN vss.gds3277
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.546 36.2835 72.606 36.4835 ;
 END
 END vss.gds3277
 PIN vss.gds3278
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 38.0475 72.774 38.2475 ;
 END
 END vss.gds3278
 PIN vss.gds3279
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.882 36.2835 72.942 36.4835 ;
 END
 END vss.gds3279
 PIN vss.gds3280
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.05 36.2835 73.11 36.4835 ;
 END
 END vss.gds3280
 PIN vss.gds3281
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.554 36.2835 73.614 36.4835 ;
 END
 END vss.gds3281
 PIN vss.gds3282
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.722 36.2835 73.782 36.4835 ;
 END
 END vss.gds3282
 PIN vss.gds3283
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.89 36.2835 73.95 36.4835 ;
 END
 END vss.gds3283
 PIN vss.gds3284
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.394 36.2835 74.454 36.4835 ;
 END
 END vss.gds3284
 PIN vss.gds3285
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.218 36.2835 73.278 36.4835 ;
 END
 END vss.gds3285
 PIN vss.gds3286
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.562 36.2835 74.622 36.4835 ;
 END
 END vss.gds3286
 PIN vss.gds3287
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.226 36.2835 74.286 36.4835 ;
 END
 END vss.gds3287
 PIN vss.gds3288
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 38.0475 70.758 38.2475 ;
 END
 END vss.gds3288
 PIN vss.gds3289
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 38.0475 73.446 38.2475 ;
 END
 END vss.gds3289
 PIN vss.gds3290
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 38.0475 74.118 38.2475 ;
 END
 END vss.gds3290
 PIN vss.gds3291
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 38.0475 74.79 38.2475 ;
 END
 END vss.gds3291
 PIN vss.gds3292
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 40.477 2.962 40.677 ;
 END
 END vss.gds3292
 PIN vss.gds3293
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 42.997 2.962 43.197 ;
 END
 END vss.gds3293
 PIN vss.gds3294
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 44.257 2.962 44.457 ;
 END
 END vss.gds3294
 PIN vss.gds3295
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 43.856 3.142 44.056 ;
 END
 END vss.gds3295
 PIN vss.gds3296
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 41.336 3.142 41.536 ;
 END
 END vss.gds3296
 PIN vss.gds3297
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 45.116 3.142 45.316 ;
 END
 END vss.gds3297
 PIN vss.gds3298
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 41.737 2.962 41.937 ;
 END
 END vss.gds3298
 PIN vss.gds3299
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 42.596 3.142 42.796 ;
 END
 END vss.gds3299
 PIN vss.gds3300
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.442 40.701 4.482 40.901 ;
 END
 END vss.gds3300
 PIN vss.gds3301
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.286 41.107 3.326 41.307 ;
 END
 END vss.gds3301
 PIN vss.gds3302
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.754 43.627 3.794 43.827 ;
 END
 END vss.gds3302
 PIN vss.gds3303
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.57 40.904 4.61 41.104 ;
 END
 END vss.gds3303
 PIN vss.gds3304
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.414 41.383 3.454 41.583 ;
 END
 END vss.gds3304
 PIN vss.gds3305
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 40.701 4.882 40.901 ;
 END
 END vss.gds3305
 PIN vss.gds3306
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 43.627 5.074 43.827 ;
 END
 END vss.gds3306
 PIN vss.gds3307
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.562 41.383 3.602 41.583 ;
 END
 END vss.gds3307
 PIN vss.gds3308
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 43.221 0.942 43.421 ;
 END
 END vss.gds3308
 PIN vss.gds3309
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 43.627 4.194 43.827 ;
 END
 END vss.gds3309
 PIN vss.gds3310
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 43.3215 0.718 43.5215 ;
 END
 END vss.gds3310
 PIN vss.gds3311
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 43.422 0.602 43.622 ;
 END
 END vss.gds3311
 PIN vss.gds3312
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 43.2305 2.122 43.4305 ;
 END
 END vss.gds3312
 PIN vss.gds3313
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 43.765 1.282 43.965 ;
 END
 END vss.gds3313
 PIN vss.gds3314
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 43.3695 1.462 43.5695 ;
 END
 END vss.gds3314
 PIN vss.gds3315
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 42.932 2.302 43.132 ;
 END
 END vss.gds3315
 PIN vss.gds3316
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 43.5235 4.002 43.7235 ;
 END
 END vss.gds3316
 PIN vss.gds3317
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 43.5235 5.282 43.7235 ;
 END
 END vss.gds3317
 PIN vss.gds3318
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 43.475 0.29 43.675 ;
 END
 END vss.gds3318
 PIN vss.gds3319
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 2.576 40.4775 2.632 40.6775 ;
 RECT 2.408 40.4775 2.464 40.6775 ;
 RECT 2.996 40.4775 3.052 40.6775 ;
 RECT 3.332 40.569 3.388 40.769 ;
 RECT 2.408 41.7375 2.464 41.9375 ;
 RECT 2.576 41.7375 2.632 41.9375 ;
 RECT 2.996 41.7375 3.052 41.9375 ;
 RECT 3.332 41.829 3.388 42.029 ;
 RECT 3.5 41.7855 3.556 41.9855 ;
 RECT 0.98 41.6525 1.036 41.8525 ;
 RECT 2.072 41.653 2.128 41.853 ;
 RECT 2.576 42.9975 2.632 43.1975 ;
 RECT 2.408 42.9975 2.464 43.1975 ;
 RECT 2.996 42.9975 3.052 43.1975 ;
 RECT 3.332 43.089 3.388 43.289 ;
 RECT 2.408 44.2575 2.464 44.4575 ;
 RECT 2.576 44.2575 2.632 44.4575 ;
 RECT 2.996 44.2575 3.052 44.4575 ;
 RECT 3.332 44.349 3.388 44.549 ;
 RECT 3.5 44.3055 3.556 44.5055 ;
 RECT 0.98 44.1725 1.036 44.3725 ;
 RECT 2.072 44.173 2.128 44.373 ;
 RECT 3.5 40.5255 3.556 40.7255 ;
 RECT 3.5 43.0455 3.556 43.2455 ;
 RECT 0.98 42.9125 1.036 43.1125 ;
 RECT 2.072 42.913 2.128 43.113 ;
 RECT 0.392 43.003 0.448 43.203 ;
 RECT 0.812 43.089 0.868 43.289 ;
 RECT 0.644 43.003 0.7 43.203 ;
 RECT 1.232 43.003 1.288 43.203 ;
 RECT 1.4 43.003 1.456 43.203 ;
 RECT 1.568 43.003 1.624 43.203 ;
 RECT 1.82 43.003 1.876 43.203 ;
 RECT 2.24 43.003 2.296 43.203 ;
 RECT 2.744 42.913 2.8 43.113 ;
 RECT 3.164 43.003 3.22 43.203 ;
 RECT 0.392 40.483 0.448 40.683 ;
 RECT 0.812 40.569 0.868 40.769 ;
 RECT 0.644 40.483 0.7 40.683 ;
 RECT 1.232 40.483 1.288 40.683 ;
 RECT 1.4 40.483 1.456 40.683 ;
 RECT 1.568 40.483 1.624 40.683 ;
 RECT 1.82 40.483 1.876 40.683 ;
 RECT 2.24 40.483 2.296 40.683 ;
 RECT 3.164 40.483 3.22 40.683 ;
 RECT 0.98 45.4325 1.036 45.6325 ;
 RECT 2.072 45.433 2.128 45.633 ;
 RECT 2.744 45.433 2.8 45.633 ;
 RECT 0.392 44.263 0.448 44.463 ;
 RECT 0.812 44.349 0.868 44.549 ;
 RECT 0.644 44.263 0.7 44.463 ;
 RECT 1.232 44.263 1.288 44.463 ;
 RECT 1.4 44.263 1.456 44.463 ;
 RECT 1.568 44.263 1.624 44.463 ;
 RECT 1.82 44.263 1.876 44.463 ;
 RECT 2.24 44.263 2.296 44.463 ;
 RECT 2.744 44.173 2.8 44.373 ;
 RECT 3.164 44.263 3.22 44.463 ;
 RECT 3.92 44.263 3.976 44.463 ;
 RECT 3.752 44.533 3.808 44.733 ;
 RECT 4.508 44.4625 4.564 44.6625 ;
 RECT 3.92 43.003 3.976 43.203 ;
 RECT 3.752 43.273 3.808 43.473 ;
 RECT 4.508 43.2025 4.564 43.4025 ;
 RECT 0.392 41.743 0.448 41.943 ;
 RECT 0.812 41.829 0.868 42.029 ;
 RECT 0.644 41.743 0.7 41.943 ;
 RECT 1.232 41.743 1.288 41.943 ;
 RECT 1.4 41.743 1.456 41.943 ;
 RECT 1.568 41.743 1.624 41.943 ;
 RECT 1.82 41.743 1.876 41.943 ;
 RECT 2.24 41.743 2.296 41.943 ;
 RECT 2.744 41.653 2.8 41.853 ;
 RECT 3.164 41.743 3.22 41.943 ;
 RECT 3.92 41.743 3.976 41.943 ;
 RECT 3.752 42.013 3.808 42.213 ;
 RECT 4.508 41.9425 4.564 42.1425 ;
 RECT 3.92 40.483 3.976 40.683 ;
 RECT 3.752 40.753 3.808 40.953 ;
 RECT 4.508 40.6825 4.564 40.8825 ;
 END
 END vss.gds3319
 PIN vss.gds3320
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.134 41.3235 10.194 41.5235 ;
 END
 END vss.gds3320
 PIN vss.gds3321
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.966 41.3235 10.026 41.5235 ;
 END
 END vss.gds3321
 PIN vss.gds3322
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.798 41.3235 9.858 41.5235 ;
 END
 END vss.gds3322
 PIN vss.gds3323
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.462 41.3235 9.522 41.5235 ;
 END
 END vss.gds3323
 PIN vss.gds3324
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.294 41.3235 9.354 41.5235 ;
 END
 END vss.gds3324
 PIN vss.gds3325
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.79 41.3235 8.85 41.5235 ;
 END
 END vss.gds3325
 PIN vss.gds3326
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.622 41.3235 8.682 41.5235 ;
 END
 END vss.gds3326
 PIN vss.gds3327
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.454 41.3235 8.514 41.5235 ;
 END
 END vss.gds3327
 PIN vss.gds3328
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.118 41.3235 8.178 41.5235 ;
 END
 END vss.gds3328
 PIN vss.gds3329
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.95 41.3235 8.01 41.5235 ;
 END
 END vss.gds3329
 PIN vss.gds3330
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.782 41.3235 7.842 41.5235 ;
 END
 END vss.gds3330
 PIN vss.gds3331
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.126 41.3235 9.186 41.5235 ;
 END
 END vss.gds3331
 PIN vss.gds3332
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.446 41.3235 7.506 41.5235 ;
 END
 END vss.gds3332
 PIN vss.gds3333
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.278 41.3235 7.338 41.5235 ;
 END
 END vss.gds3333
 PIN vss.gds3334
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 42.9595 9.69 43.1595 ;
 END
 END vss.gds3334
 PIN vss.gds3335
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 42.9595 9.018 43.1595 ;
 END
 END vss.gds3335
 PIN vss.gds3336
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.11 41.3235 7.17 41.5235 ;
 END
 END vss.gds3336
 PIN vss.gds3337
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 43.424 6.178 43.624 ;
 END
 END vss.gds3337
 PIN vss.gds3338
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 43.627 5.474 43.827 ;
 END
 END vss.gds3338
 PIN vss.gds3339
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 42.9595 8.346 43.1595 ;
 END
 END vss.gds3339
 PIN vss.gds3340
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 42.9595 7.674 43.1595 ;
 END
 END vss.gds3340
 PIN vss.gds3341
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 43.627 5.73 43.827 ;
 END
 END vss.gds3341
 PIN vss.gds3342
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 43.627 5.986 43.827 ;
 END
 END vss.gds3342
 PIN vss.gds3343
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 43.233 6.434 43.433 ;
 END
 END vss.gds3343
 PIN vss.gds3344
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 6.608 44.533 6.664 44.733 ;
 RECT 6.524 44.256 6.58 44.456 ;
 RECT 6.692 44.406 6.748 44.606 ;
 RECT 6.692 43.146 6.748 43.346 ;
 RECT 6.524 42.996 6.58 43.196 ;
 RECT 6.608 43.273 6.664 43.473 ;
 RECT 6.608 42.013 6.664 42.213 ;
 RECT 6.524 41.736 6.58 41.936 ;
 RECT 6.692 41.886 6.748 42.086 ;
 RECT 6.692 40.626 6.748 40.826 ;
 RECT 6.524 40.476 6.58 40.676 ;
 RECT 6.608 40.753 6.664 40.953 ;
 END
 END vss.gds3344
 PIN vss.gds3345
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 42.242 13.898 42.442 ;
 END
 END vss.gds3345
 PIN vss.gds3346
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 42.282 14.87 42.482 ;
 END
 END vss.gds3346
 PIN vss.gds3347
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 40.982 13.898 41.182 ;
 END
 END vss.gds3347
 PIN vss.gds3348
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 41.022 14.87 41.222 ;
 END
 END vss.gds3348
 PIN vss.gds3349
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 43.502 13.898 43.702 ;
 END
 END vss.gds3349
 PIN vss.gds3350
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 43.542 14.87 43.742 ;
 END
 END vss.gds3350
 PIN vss.gds3351
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 44.762 13.898 44.962 ;
 END
 END vss.gds3351
 PIN vss.gds3352
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 44.802 14.87 45.002 ;
 END
 END vss.gds3352
 PIN vss.gds3353
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.15 41.3235 12.21 41.5235 ;
 END
 END vss.gds3353
 PIN vss.gds3354
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.982 41.3235 12.042 41.5235 ;
 END
 END vss.gds3354
 PIN vss.gds3355
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.814 41.3235 11.874 41.5235 ;
 END
 END vss.gds3355
 PIN vss.gds3356
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.478 41.3235 11.538 41.5235 ;
 END
 END vss.gds3356
 PIN vss.gds3357
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.31 41.3235 11.37 41.5235 ;
 END
 END vss.gds3357
 PIN vss.gds3358
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.142 41.3235 11.202 41.5235 ;
 END
 END vss.gds3358
 PIN vss.gds3359
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.806 41.3235 10.866 41.5235 ;
 END
 END vss.gds3359
 PIN vss.gds3360
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.638 41.3235 10.698 41.5235 ;
 END
 END vss.gds3360
 PIN vss.gds3361
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.47 41.3235 10.53 41.5235 ;
 END
 END vss.gds3361
 PIN vss.gds3362
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 42.0095 13.058 42.2095 ;
 END
 END vss.gds3362
 PIN vss.gds3363
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.262 44.316 13.318 44.516 ;
 END
 END vss.gds3363
 PIN vss.gds3364
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 42.9595 11.706 43.1595 ;
 END
 END vss.gds3364
 PIN vss.gds3365
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 42.9595 11.034 43.1595 ;
 END
 END vss.gds3365
 PIN vss.gds3366
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 42.9595 10.362 43.1595 ;
 END
 END vss.gds3366
 PIN vss.gds3367
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 43.128 15.162 43.328 ;
 END
 END vss.gds3367
 PIN vss.gds3368
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 43.128 14.498 43.328 ;
 END
 END vss.gds3368
 PIN vss.gds3369
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 42.9595 13.658 43.1595 ;
 END
 END vss.gds3369
 PIN vss.gds3370
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 42.925 12.378 43.125 ;
 END
 END vss.gds3370
 PIN vss.gds3371
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 43.627 12.59 43.827 ;
 END
 END vss.gds3371
 PIN vss.gds3372
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 43.1235 12.818 43.3235 ;
 END
 END vss.gds3372
 PIN vss.gds3373
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 14 44.94 14.056 45.113 ;
 RECT 14.168 44.913 14.224 45.113 ;
 RECT 14 43.68 14.056 43.853 ;
 RECT 14.168 43.653 14.224 43.853 ;
 RECT 14 41.16 14.056 41.333 ;
 RECT 14.168 41.133 14.224 41.333 ;
 RECT 14 42.42 14.056 42.593 ;
 RECT 14.168 42.393 14.224 42.593 ;
 RECT 14.336 41.753 14.392 41.953 ;
 RECT 14.168 41.753 14.224 41.953 ;
 RECT 14.336 40.493 14.392 40.693 ;
 RECT 14.168 40.493 14.224 40.693 ;
 RECT 14.336 43.013 14.392 43.213 ;
 RECT 14.168 43.013 14.224 43.213 ;
 RECT 14.336 44.273 14.392 44.473 ;
 RECT 14.168 44.273 14.224 44.473 ;
 RECT 13.664 41.887 13.72 42.087 ;
 RECT 15.008 41.963 15.064 42.163 ;
 RECT 14.84 42.437 14.896 42.602 ;
 RECT 14.672 42.437 14.728 42.602 ;
 RECT 13.664 40.627 13.72 40.827 ;
 RECT 15.008 40.703 15.064 40.903 ;
 RECT 14.84 41.177 14.896 41.342 ;
 RECT 14.672 41.177 14.728 41.342 ;
 RECT 15.008 43.223 15.064 43.423 ;
 RECT 14.84 43.697 14.896 43.862 ;
 RECT 14.672 43.697 14.728 43.862 ;
 RECT 13.664 43.147 13.72 43.347 ;
 RECT 15.008 44.483 15.064 44.683 ;
 RECT 14.84 44.957 14.896 45.122 ;
 RECT 14.672 44.957 14.728 45.122 ;
 RECT 13.664 44.407 13.72 44.607 ;
 RECT 15.176 41.4035 15.232 41.6035 ;
 RECT 12.824 41.188 12.88 41.388 ;
 RECT 13.496 41.199 13.552 41.399 ;
 RECT 13.328 41.137 13.384 41.337 ;
 RECT 13.16 41.188 13.216 41.388 ;
 RECT 12.488 41.218 12.544 41.418 ;
 RECT 12.992 41.188 13.048 41.388 ;
 RECT 12.656 41.218 12.712 41.418 ;
 END
 END vss.gds3373
 PIN vss.gds3374
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 40.477 16.146 40.677 ;
 END
 END vss.gds3374
 PIN vss.gds3375
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 45 15.418 45.2 ;
 END
 END vss.gds3375
 PIN vss.gds3376
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.438 43.8995 17.494 44.0995 ;
 END
 END vss.gds3376
 PIN vss.gds3377
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 42.9595 20.274 43.1595 ;
 END
 END vss.gds3377
 PIN vss.gds3378
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.702 41.3235 18.762 41.5235 ;
 END
 END vss.gds3378
 PIN vss.gds3379
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 44.257 16.146 44.457 ;
 END
 END vss.gds3379
 PIN vss.gds3380
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 42.997 16.146 43.197 ;
 END
 END vss.gds3380
 PIN vss.gds3381
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 41.737 16.146 41.937 ;
 END
 END vss.gds3381
 PIN vss.gds3382
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.038 41.3235 19.098 41.5235 ;
 END
 END vss.gds3382
 PIN vss.gds3383
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.206 41.3235 19.266 41.5235 ;
 END
 END vss.gds3383
 PIN vss.gds3384
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.374 41.3235 19.434 41.5235 ;
 END
 END vss.gds3384
 PIN vss.gds3385
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.71 41.3235 19.77 41.5235 ;
 END
 END vss.gds3385
 PIN vss.gds3386
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.878 41.3235 19.938 41.5235 ;
 END
 END vss.gds3386
 PIN vss.gds3387
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.534 41.3235 18.594 41.5235 ;
 END
 END vss.gds3387
 PIN vss.gds3388
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 41.796 16.814 41.996 ;
 END
 END vss.gds3388
 PIN vss.gds3389
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.366 41.3235 18.426 41.5235 ;
 END
 END vss.gds3389
 PIN vss.gds3390
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 44.7555 17.314 44.9555 ;
 END
 END vss.gds3390
 PIN vss.gds3391
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.986 41.107 18.026 41.307 ;
 END
 END vss.gds3391
 PIN vss.gds3392
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 42.9595 18.93 43.1595 ;
 END
 END vss.gds3392
 PIN vss.gds3393
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 42.9595 19.602 43.1595 ;
 END
 END vss.gds3393
 PIN vss.gds3394
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 43.0465 16.994 43.2465 ;
 END
 END vss.gds3394
 PIN vss.gds3395
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.046 41.3235 20.106 41.5235 ;
 END
 END vss.gds3395
 PIN vss.gds3396
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 43.128 15.842 43.328 ;
 END
 END vss.gds3396
 PIN vss.gds3397
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 42.925 18.258 43.125 ;
 END
 END vss.gds3397
 PIN vss.gds3398
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 43.1235 17.834 43.3235 ;
 END
 END vss.gds3398
 PIN vss.gds3399
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 43.2305 16.49 43.4305 ;
 END
 END vss.gds3399
 PIN vss.gds3400
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 15.596 45.184 15.652 45.384 ;
 RECT 15.848 45.187 15.904 45.387 ;
 RECT 15.596 43.924 15.652 44.124 ;
 RECT 15.848 43.927 15.904 44.127 ;
 RECT 16.52 44.96 16.576 45.113 ;
 RECT 15.764 44.957 15.82 45.122 ;
 RECT 15.596 44.957 15.652 45.122 ;
 RECT 15.596 42.664 15.652 42.864 ;
 RECT 15.848 42.667 15.904 42.867 ;
 RECT 16.52 43.7 16.576 43.853 ;
 RECT 15.764 43.697 15.82 43.862 ;
 RECT 15.596 43.697 15.652 43.862 ;
 RECT 16.52 41.18 16.576 41.333 ;
 RECT 15.764 41.177 15.82 41.342 ;
 RECT 15.596 41.177 15.652 41.342 ;
 RECT 15.596 41.404 15.652 41.604 ;
 RECT 15.848 41.407 15.904 41.607 ;
 RECT 16.52 42.44 16.576 42.593 ;
 RECT 15.764 42.437 15.82 42.602 ;
 RECT 15.596 42.437 15.652 42.602 ;
 RECT 16.856 40.5515 16.912 40.7515 ;
 RECT 16.352 40.8035 16.408 41.0035 ;
 RECT 16.352 42.0635 16.408 42.2635 ;
 RECT 16.856 41.8115 16.912 42.0115 ;
 RECT 15.428 41.963 15.484 42.163 ;
 RECT 15.428 40.703 15.484 40.903 ;
 RECT 15.428 43.223 15.484 43.423 ;
 RECT 16.352 43.3235 16.408 43.5235 ;
 RECT 16.856 43.0715 16.912 43.2715 ;
 RECT 15.428 44.483 15.484 44.683 ;
 RECT 16.352 44.5835 16.408 44.7835 ;
 RECT 16.856 44.3315 16.912 44.5315 ;
 RECT 17.864 41.218 17.92 41.418 ;
 RECT 17.696 41.2255 17.752 41.4255 ;
 RECT 17.528 41.218 17.584 41.418 ;
 RECT 17.36 41.218 17.416 41.418 ;
 RECT 17.192 41.218 17.248 41.418 ;
 RECT 18.032 41.218 18.088 41.418 ;
 RECT 17.024 41.333 17.08 41.533 ;
 END
 END vss.gds3400
 PIN vss.gds3401
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.17 41.3235 25.23 41.5235 ;
 END
 END vss.gds3401
 PIN vss.gds3402
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.002 41.3235 25.062 41.5235 ;
 END
 END vss.gds3402
 PIN vss.gds3403
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.834 41.3235 24.894 41.5235 ;
 END
 END vss.gds3403
 PIN vss.gds3404
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.498 41.3235 24.558 41.5235 ;
 END
 END vss.gds3404
 PIN vss.gds3405
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.33 41.3235 24.39 41.5235 ;
 END
 END vss.gds3405
 PIN vss.gds3406
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.162 41.3235 24.222 41.5235 ;
 END
 END vss.gds3406
 PIN vss.gds3407
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.382 41.3235 20.442 41.5235 ;
 END
 END vss.gds3407
 PIN vss.gds3408
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.55 41.3235 20.61 41.5235 ;
 END
 END vss.gds3408
 PIN vss.gds3409
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.718 41.3235 20.778 41.5235 ;
 END
 END vss.gds3409
 PIN vss.gds3410
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.054 41.3235 21.114 41.5235 ;
 END
 END vss.gds3410
 PIN vss.gds3411
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.222 41.3235 21.282 41.5235 ;
 END
 END vss.gds3411
 PIN vss.gds3412
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.39 41.3235 21.45 41.5235 ;
 END
 END vss.gds3412
 PIN vss.gds3413
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.726 41.3235 21.786 41.5235 ;
 END
 END vss.gds3413
 PIN vss.gds3414
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.894 41.3235 21.954 41.5235 ;
 END
 END vss.gds3414
 PIN vss.gds3415
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.062 41.3235 22.122 41.5235 ;
 END
 END vss.gds3415
 PIN vss.gds3416
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 42.9595 24.726 43.1595 ;
 END
 END vss.gds3416
 PIN vss.gds3417
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 42.9595 21.618 43.1595 ;
 END
 END vss.gds3417
 PIN vss.gds3418
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 42.9595 20.946 43.1595 ;
 END
 END vss.gds3418
 PIN vss.gds3419
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 42.9595 22.29 43.1595 ;
 END
 END vss.gds3419
 PIN vss.gds3420
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.398 41.3235 22.458 41.5235 ;
 END
 END vss.gds3420
 PIN vss.gds3421
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.566 41.3235 22.626 41.5235 ;
 END
 END vss.gds3421
 PIN vss.gds3422
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.734 41.3235 22.794 41.5235 ;
 END
 END vss.gds3422
 PIN vss.gds3423
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.07 41.3235 23.13 41.5235 ;
 END
 END vss.gds3423
 PIN vss.gds3424
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.238 41.3235 23.298 41.5235 ;
 END
 END vss.gds3424
 PIN vss.gds3425
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.406 41.3235 23.466 41.5235 ;
 END
 END vss.gds3425
 PIN vss.gds3426
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 42.9595 22.962 43.1595 ;
 END
 END vss.gds3426
 PIN vss.gds3427
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 42.9595 23.634 43.1595 ;
 END
 END vss.gds3427
 PIN vss.gds3428
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 23.912 40.64 23.968 40.84 ;
 RECT 23.912 41.9 23.968 42.1 ;
 RECT 23.912 43.16 23.968 43.36 ;
 RECT 23.912 44.42 23.968 44.62 ;
 RECT 23.744 43.09 23.8 43.29 ;
 END
 END vss.gds3428
 PIN vss.gds3429
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.202 41.3235 29.262 41.5235 ;
 END
 END vss.gds3429
 PIN vss.gds3430
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.034 41.3235 29.094 41.5235 ;
 END
 END vss.gds3430
 PIN vss.gds3431
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.866 41.3235 28.926 41.5235 ;
 END
 END vss.gds3431
 PIN vss.gds3432
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.53 41.3235 28.59 41.5235 ;
 END
 END vss.gds3432
 PIN vss.gds3433
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.362 41.3235 28.422 41.5235 ;
 END
 END vss.gds3433
 PIN vss.gds3434
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.194 41.3235 28.254 41.5235 ;
 END
 END vss.gds3434
 PIN vss.gds3435
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.858 41.3235 27.918 41.5235 ;
 END
 END vss.gds3435
 PIN vss.gds3436
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.69 41.3235 27.75 41.5235 ;
 END
 END vss.gds3436
 PIN vss.gds3437
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.522 41.3235 27.582 41.5235 ;
 END
 END vss.gds3437
 PIN vss.gds3438
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.186 41.3235 27.246 41.5235 ;
 END
 END vss.gds3438
 PIN vss.gds3439
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.018 41.3235 27.078 41.5235 ;
 END
 END vss.gds3439
 PIN vss.gds3440
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.85 41.3235 26.91 41.5235 ;
 END
 END vss.gds3440
 PIN vss.gds3441
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.514 41.3235 26.574 41.5235 ;
 END
 END vss.gds3441
 PIN vss.gds3442
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.346 41.3235 26.406 41.5235 ;
 END
 END vss.gds3442
 PIN vss.gds3443
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.178 41.3235 26.238 41.5235 ;
 END
 END vss.gds3443
 PIN vss.gds3444
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.842 41.3235 25.902 41.5235 ;
 END
 END vss.gds3444
 PIN vss.gds3445
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.674 41.3235 25.734 41.5235 ;
 END
 END vss.gds3445
 PIN vss.gds3446
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.506 41.3235 25.566 41.5235 ;
 END
 END vss.gds3446
 PIN vss.gds3447
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 42.9595 28.758 43.1595 ;
 END
 END vss.gds3447
 PIN vss.gds3448
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 42.9595 28.086 43.1595 ;
 END
 END vss.gds3448
 PIN vss.gds3449
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 42.9595 27.414 43.1595 ;
 END
 END vss.gds3449
 PIN vss.gds3450
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 42.9595 26.742 43.1595 ;
 END
 END vss.gds3450
 PIN vss.gds3451
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 42.9595 26.07 43.1595 ;
 END
 END vss.gds3451
 PIN vss.gds3452
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 42.9595 25.398 43.1595 ;
 END
 END vss.gds3452
 PIN vss.gds3453
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 42.925 29.43 43.125 ;
 END
 END vss.gds3453
 PIN vss.gds3454
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 42.0095 30.11 42.2095 ;
 END
 END vss.gds3454
 PIN vss.gds3455
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 43.1235 29.87 43.3235 ;
 END
 END vss.gds3455
 PIN vss.gds3456
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 43.627 29.642 43.827 ;
 END
 END vss.gds3456
 PIN vss.gds3457
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.876 41.188 29.932 41.388 ;
 RECT 29.708 41.218 29.764 41.418 ;
 RECT 30.212 41.188 30.268 41.388 ;
 RECT 29.54 41.218 29.596 41.418 ;
 RECT 30.044 41.188 30.1 41.388 ;
 END
 END vss.gds3457
 PIN vss.gds3458
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 42.282 31.922 42.482 ;
 END
 END vss.gds3458
 PIN vss.gds3459
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 41.022 31.922 41.222 ;
 END
 END vss.gds3459
 PIN vss.gds3460
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 43.542 31.922 43.742 ;
 END
 END vss.gds3460
 PIN vss.gds3461
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 44.802 31.922 45.002 ;
 END
 END vss.gds3461
 PIN vss.gds3462
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 40.982 30.95 41.182 ;
 END
 END vss.gds3462
 PIN vss.gds3463
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.314 44.316 30.37 44.516 ;
 END
 END vss.gds3463
 PIN vss.gds3464
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 44.762 30.95 44.962 ;
 END
 END vss.gds3464
 PIN vss.gds3465
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 44.257 33.198 44.457 ;
 END
 END vss.gds3465
 PIN vss.gds3466
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 42.997 33.198 43.197 ;
 END
 END vss.gds3466
 PIN vss.gds3467
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.49 43.8995 34.546 44.0995 ;
 END
 END vss.gds3467
 PIN vss.gds3468
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 41.737 33.198 41.937 ;
 END
 END vss.gds3468
 PIN vss.gds3469
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 40.477 33.198 40.677 ;
 END
 END vss.gds3469
 PIN vss.gds3470
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 41.796 33.866 41.996 ;
 END
 END vss.gds3470
 PIN vss.gds3471
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 43.128 32.214 43.328 ;
 END
 END vss.gds3471
 PIN vss.gds3472
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 43.0465 34.046 43.2465 ;
 END
 END vss.gds3472
 PIN vss.gds3473
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 43.502 30.95 43.702 ;
 END
 END vss.gds3473
 PIN vss.gds3474
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 42.242 30.95 42.442 ;
 END
 END vss.gds3474
 PIN vss.gds3475
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 44.7555 34.366 44.9555 ;
 END
 END vss.gds3475
 PIN vss.gds3476
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 45 32.47 45.2 ;
 END
 END vss.gds3476
 PIN vss.gds3477
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.038 41.107 35.078 41.307 ;
 END
 END vss.gds3477
 PIN vss.gds3478
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 42.9595 30.71 43.1595 ;
 END
 END vss.gds3478
 PIN vss.gds3479
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 43.128 32.894 43.328 ;
 END
 END vss.gds3479
 PIN vss.gds3480
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 43.2305 33.542 43.4305 ;
 END
 END vss.gds3480
 PIN vss.gds3481
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 43.128 31.55 43.328 ;
 END
 END vss.gds3481
 PIN vss.gds3482
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 43.1235 34.886 43.3235 ;
 END
 END vss.gds3482
 PIN vss.gds3483
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 32.648 45.184 32.704 45.384 ;
 RECT 32.9 45.187 32.956 45.387 ;
 RECT 32.648 43.924 32.704 44.124 ;
 RECT 32.9 43.927 32.956 44.127 ;
 RECT 33.572 44.96 33.628 45.113 ;
 RECT 31.052 44.94 31.108 45.113 ;
 RECT 31.22 44.913 31.276 45.113 ;
 RECT 32.816 44.957 32.872 45.122 ;
 RECT 32.648 44.957 32.704 45.122 ;
 RECT 31.892 44.957 31.948 45.122 ;
 RECT 31.724 44.957 31.78 45.122 ;
 RECT 32.648 42.664 32.704 42.864 ;
 RECT 32.9 42.667 32.956 42.867 ;
 RECT 33.572 43.7 33.628 43.853 ;
 RECT 31.052 43.68 31.108 43.853 ;
 RECT 31.22 43.653 31.276 43.853 ;
 RECT 32.816 43.697 32.872 43.862 ;
 RECT 32.648 43.697 32.704 43.862 ;
 RECT 31.892 43.697 31.948 43.862 ;
 RECT 31.724 43.697 31.78 43.862 ;
 RECT 33.572 41.18 33.628 41.333 ;
 RECT 31.052 41.16 31.108 41.333 ;
 RECT 31.22 41.133 31.276 41.333 ;
 RECT 32.816 41.177 32.872 41.342 ;
 RECT 32.648 41.177 32.704 41.342 ;
 RECT 31.892 41.177 31.948 41.342 ;
 RECT 31.724 41.177 31.78 41.342 ;
 RECT 33.572 42.44 33.628 42.593 ;
 RECT 31.052 42.42 31.108 42.593 ;
 RECT 31.22 42.393 31.276 42.593 ;
 RECT 32.816 42.437 32.872 42.602 ;
 RECT 32.648 42.437 32.704 42.602 ;
 RECT 31.892 42.437 31.948 42.602 ;
 RECT 31.724 42.437 31.78 42.602 ;
 RECT 32.648 41.404 32.704 41.604 ;
 RECT 32.9 41.407 32.956 41.607 ;
 RECT 32.06 44.483 32.116 44.683 ;
 RECT 31.388 44.273 31.444 44.473 ;
 RECT 31.22 44.273 31.276 44.473 ;
 RECT 32.48 44.483 32.536 44.683 ;
 RECT 31.388 43.013 31.444 43.213 ;
 RECT 31.22 43.013 31.276 43.213 ;
 RECT 32.06 43.223 32.116 43.423 ;
 RECT 32.48 43.223 32.536 43.423 ;
 RECT 31.388 41.753 31.444 41.953 ;
 RECT 31.22 41.753 31.276 41.953 ;
 RECT 32.06 41.963 32.116 42.163 ;
 RECT 32.48 41.963 32.536 42.163 ;
 RECT 33.908 40.5515 33.964 40.7515 ;
 RECT 33.404 40.8035 33.46 41.0035 ;
 RECT 32.06 40.703 32.116 40.903 ;
 RECT 32.48 40.703 32.536 40.903 ;
 RECT 31.388 40.493 31.444 40.693 ;
 RECT 31.22 40.493 31.276 40.693 ;
 RECT 30.716 40.627 30.772 40.827 ;
 RECT 30.716 41.887 30.772 42.087 ;
 RECT 33.404 42.0635 33.46 42.2635 ;
 RECT 33.908 41.8115 33.964 42.0115 ;
 RECT 30.716 43.147 30.772 43.347 ;
 RECT 33.404 43.3235 33.46 43.5235 ;
 RECT 33.908 43.0715 33.964 43.2715 ;
 RECT 30.716 44.407 30.772 44.607 ;
 RECT 33.404 44.5835 33.46 44.7835 ;
 RECT 33.908 44.3315 33.964 44.5315 ;
 RECT 30.548 41.199 30.604 41.399 ;
 RECT 34.916 41.218 34.972 41.418 ;
 RECT 32.228 41.4035 32.284 41.6035 ;
 RECT 30.38 41.137 30.436 41.337 ;
 RECT 34.748 41.2255 34.804 41.4255 ;
 RECT 34.58 41.218 34.636 41.418 ;
 RECT 34.412 41.218 34.468 41.418 ;
 RECT 34.244 41.218 34.3 41.418 ;
 RECT 34.076 41.333 34.132 41.533 ;
 RECT 35.084 41.218 35.14 41.418 ;
 END
 END vss.gds3483
 PIN vss.gds3484
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.122 41.3235 40.182 41.5235 ;
 END
 END vss.gds3484
 PIN vss.gds3485
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.754 41.3235 35.814 41.5235 ;
 END
 END vss.gds3485
 PIN vss.gds3486
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.09 41.3235 36.15 41.5235 ;
 END
 END vss.gds3486
 PIN vss.gds3487
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.258 41.3235 36.318 41.5235 ;
 END
 END vss.gds3487
 PIN vss.gds3488
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.426 41.3235 36.486 41.5235 ;
 END
 END vss.gds3488
 PIN vss.gds3489
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 42.9595 36.654 43.1595 ;
 END
 END vss.gds3489
 PIN vss.gds3490
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.762 41.3235 36.822 41.5235 ;
 END
 END vss.gds3490
 PIN vss.gds3491
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.93 41.3235 36.99 41.5235 ;
 END
 END vss.gds3491
 PIN vss.gds3492
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.098 41.3235 37.158 41.5235 ;
 END
 END vss.gds3492
 PIN vss.gds3493
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 42.9595 37.326 43.1595 ;
 END
 END vss.gds3493
 PIN vss.gds3494
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.434 41.3235 37.494 41.5235 ;
 END
 END vss.gds3494
 PIN vss.gds3495
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.602 41.3235 37.662 41.5235 ;
 END
 END vss.gds3495
 PIN vss.gds3496
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.77 41.3235 37.83 41.5235 ;
 END
 END vss.gds3496
 PIN vss.gds3497
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 42.9595 37.998 43.1595 ;
 END
 END vss.gds3497
 PIN vss.gds3498
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.106 41.3235 38.166 41.5235 ;
 END
 END vss.gds3498
 PIN vss.gds3499
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.274 41.3235 38.334 41.5235 ;
 END
 END vss.gds3499
 PIN vss.gds3500
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.442 41.3235 38.502 41.5235 ;
 END
 END vss.gds3500
 PIN vss.gds3501
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.778 41.3235 38.838 41.5235 ;
 END
 END vss.gds3501
 PIN vss.gds3502
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.946 41.3235 39.006 41.5235 ;
 END
 END vss.gds3502
 PIN vss.gds3503
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.45 41.3235 39.51 41.5235 ;
 END
 END vss.gds3503
 PIN vss.gds3504
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.618 41.3235 39.678 41.5235 ;
 END
 END vss.gds3504
 PIN vss.gds3505
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.586 41.3235 35.646 41.5235 ;
 END
 END vss.gds3505
 PIN vss.gds3506
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.786 41.3235 39.846 41.5235 ;
 END
 END vss.gds3506
 PIN vss.gds3507
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.114 41.3235 39.174 41.5235 ;
 END
 END vss.gds3507
 PIN vss.gds3508
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.418 41.3235 35.478 41.5235 ;
 END
 END vss.gds3508
 PIN vss.gds3509
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 42.9595 38.67 43.1595 ;
 END
 END vss.gds3509
 PIN vss.gds3510
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 42.9595 35.982 43.1595 ;
 END
 END vss.gds3510
 PIN vss.gds3511
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 42.9595 40.014 43.1595 ;
 END
 END vss.gds3511
 PIN vss.gds3512
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 42.925 35.31 43.125 ;
 END
 END vss.gds3512
 PIN vss.gds3513
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 42.9595 39.342 43.1595 ;
 END
 END vss.gds3513
 PIN vss.gds3514
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 42.9595 45.138 43.1595 ;
 END
 END vss.gds3514
 PIN vss.gds3515
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.91 41.3235 44.97 41.5235 ;
 END
 END vss.gds3515
 PIN vss.gds3516
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.742 41.3235 44.802 41.5235 ;
 END
 END vss.gds3516
 PIN vss.gds3517
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.574 41.3235 44.634 41.5235 ;
 END
 END vss.gds3517
 PIN vss.gds3518
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 42.9595 44.466 43.1595 ;
 END
 END vss.gds3518
 PIN vss.gds3519
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.238 41.3235 44.298 41.5235 ;
 END
 END vss.gds3519
 PIN vss.gds3520
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.07 41.3235 44.13 41.5235 ;
 END
 END vss.gds3520
 PIN vss.gds3521
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.902 41.3235 43.962 41.5235 ;
 END
 END vss.gds3521
 PIN vss.gds3522
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 42.9595 43.794 43.1595 ;
 END
 END vss.gds3522
 PIN vss.gds3523
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.566 41.3235 43.626 41.5235 ;
 END
 END vss.gds3523
 PIN vss.gds3524
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.398 41.3235 43.458 41.5235 ;
 END
 END vss.gds3524
 PIN vss.gds3525
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.23 41.3235 43.29 41.5235 ;
 END
 END vss.gds3525
 PIN vss.gds3526
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 42.9595 43.122 43.1595 ;
 END
 END vss.gds3526
 PIN vss.gds3527
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.894 41.3235 42.954 41.5235 ;
 END
 END vss.gds3527
 PIN vss.gds3528
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.726 41.3235 42.786 41.5235 ;
 END
 END vss.gds3528
 PIN vss.gds3529
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.558 41.3235 42.618 41.5235 ;
 END
 END vss.gds3529
 PIN vss.gds3530
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 42.9595 42.45 43.1595 ;
 END
 END vss.gds3530
 PIN vss.gds3531
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.222 41.3235 42.282 41.5235 ;
 END
 END vss.gds3531
 PIN vss.gds3532
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.054 41.3235 42.114 41.5235 ;
 END
 END vss.gds3532
 PIN vss.gds3533
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.886 41.3235 41.946 41.5235 ;
 END
 END vss.gds3533
 PIN vss.gds3534
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 42.9595 41.778 43.1595 ;
 END
 END vss.gds3534
 PIN vss.gds3535
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.55 41.3235 41.61 41.5235 ;
 END
 END vss.gds3535
 PIN vss.gds3536
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.382 41.3235 41.442 41.5235 ;
 END
 END vss.gds3536
 PIN vss.gds3537
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.214 41.3235 41.274 41.5235 ;
 END
 END vss.gds3537
 PIN vss.gds3538
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.29 41.3235 40.35 41.5235 ;
 END
 END vss.gds3538
 PIN vss.gds3539
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.458 41.3235 40.518 41.5235 ;
 END
 END vss.gds3539
 PIN vss.gds3540
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 42.9595 40.686 43.1595 ;
 END
 END vss.gds3540
 PIN vss.gds3541
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 40.964 44.42 41.02 44.62 ;
 RECT 40.964 43.16 41.02 43.36 ;
 RECT 40.964 41.9 41.02 42.1 ;
 RECT 40.964 40.64 41.02 40.84 ;
 RECT 40.796 43.09 40.852 43.29 ;
 END
 END vss.gds3541
 PIN vss.gds3542
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 42.282 48.974 42.482 ;
 END
 END vss.gds3542
 PIN vss.gds3543
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 41.022 48.974 41.222 ;
 END
 END vss.gds3543
 PIN vss.gds3544
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 43.542 48.974 43.742 ;
 END
 END vss.gds3544
 PIN vss.gds3545
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 44.802 48.974 45.002 ;
 END
 END vss.gds3545
 PIN vss.gds3546
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 40.982 48.002 41.182 ;
 END
 END vss.gds3546
 PIN vss.gds3547
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 43.502 48.002 43.702 ;
 END
 END vss.gds3547
 PIN vss.gds3548
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 44.762 48.002 44.962 ;
 END
 END vss.gds3548
 PIN vss.gds3549
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.366 44.316 47.422 44.516 ;
 END
 END vss.gds3549
 PIN vss.gds3550
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 42.925 46.482 43.125 ;
 END
 END vss.gds3550
 PIN vss.gds3551
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.254 41.3235 46.314 41.5235 ;
 END
 END vss.gds3551
 PIN vss.gds3552
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.086 41.3235 46.146 41.5235 ;
 END
 END vss.gds3552
 PIN vss.gds3553
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.918 41.3235 45.978 41.5235 ;
 END
 END vss.gds3553
 PIN vss.gds3554
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 42.9595 45.81 43.1595 ;
 END
 END vss.gds3554
 PIN vss.gds3555
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.582 41.3235 45.642 41.5235 ;
 END
 END vss.gds3555
 PIN vss.gds3556
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.414 41.3235 45.474 41.5235 ;
 END
 END vss.gds3556
 PIN vss.gds3557
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.246 41.3235 45.306 41.5235 ;
 END
 END vss.gds3557
 PIN vss.gds3558
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 44.257 50.25 44.457 ;
 END
 END vss.gds3558
 PIN vss.gds3559
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 42.997 50.25 43.197 ;
 END
 END vss.gds3559
 PIN vss.gds3560
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 42.0095 47.162 42.2095 ;
 END
 END vss.gds3560
 PIN vss.gds3561
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 45 49.522 45.2 ;
 END
 END vss.gds3561
 PIN vss.gds3562
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 41.737 50.25 41.937 ;
 END
 END vss.gds3562
 PIN vss.gds3563
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 42.242 48.002 42.442 ;
 END
 END vss.gds3563
 PIN vss.gds3564
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 40.477 50.25 40.677 ;
 END
 END vss.gds3564
 PIN vss.gds3565
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 43.1235 46.922 43.3235 ;
 END
 END vss.gds3565
 PIN vss.gds3566
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 43.627 46.694 43.827 ;
 END
 END vss.gds3566
 PIN vss.gds3567
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 42.9595 47.762 43.1595 ;
 END
 END vss.gds3567
 PIN vss.gds3568
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 43.128 49.266 43.328 ;
 END
 END vss.gds3568
 PIN vss.gds3569
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 43.128 48.602 43.328 ;
 END
 END vss.gds3569
 PIN vss.gds3570
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 43.128 49.946 43.328 ;
 END
 END vss.gds3570
 PIN vss.gds3571
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 49.7 43.924 49.756 44.124 ;
 RECT 49.952 43.927 50.008 44.127 ;
 RECT 48.104 44.94 48.16 45.113 ;
 RECT 48.272 44.913 48.328 45.113 ;
 RECT 49.868 44.957 49.924 45.122 ;
 RECT 49.7 44.957 49.756 45.122 ;
 RECT 48.944 44.957 49 45.122 ;
 RECT 48.776 44.957 48.832 45.122 ;
 RECT 49.7 42.664 49.756 42.864 ;
 RECT 49.952 42.667 50.008 42.867 ;
 RECT 48.104 43.68 48.16 43.853 ;
 RECT 48.272 43.653 48.328 43.853 ;
 RECT 49.868 43.697 49.924 43.862 ;
 RECT 49.7 43.697 49.756 43.862 ;
 RECT 48.944 43.697 49 43.862 ;
 RECT 48.776 43.697 48.832 43.862 ;
 RECT 48.104 41.16 48.16 41.333 ;
 RECT 48.272 41.133 48.328 41.333 ;
 RECT 49.868 41.177 49.924 41.342 ;
 RECT 49.7 41.177 49.756 41.342 ;
 RECT 48.944 41.177 49 41.342 ;
 RECT 48.776 41.177 48.832 41.342 ;
 RECT 48.104 42.42 48.16 42.593 ;
 RECT 48.272 42.393 48.328 42.593 ;
 RECT 49.868 42.437 49.924 42.602 ;
 RECT 49.7 42.437 49.756 42.602 ;
 RECT 48.944 42.437 49 42.602 ;
 RECT 48.776 42.437 48.832 42.602 ;
 RECT 49.7 41.404 49.756 41.604 ;
 RECT 49.952 41.407 50.008 41.607 ;
 RECT 49.7 45.184 49.756 45.384 ;
 RECT 49.952 45.187 50.008 45.387 ;
 RECT 49.112 44.483 49.168 44.683 ;
 RECT 48.44 44.273 48.496 44.473 ;
 RECT 48.272 44.273 48.328 44.473 ;
 RECT 47.768 44.407 47.824 44.607 ;
 RECT 49.532 44.483 49.588 44.683 ;
 RECT 48.44 41.753 48.496 41.953 ;
 RECT 48.272 41.753 48.328 41.953 ;
 RECT 49.112 41.963 49.168 42.163 ;
 RECT 49.532 41.963 49.588 42.163 ;
 RECT 49.112 40.703 49.168 40.903 ;
 RECT 48.44 40.493 48.496 40.693 ;
 RECT 48.272 40.493 48.328 40.693 ;
 RECT 49.112 43.223 49.168 43.423 ;
 RECT 49.532 43.223 49.588 43.423 ;
 RECT 48.44 43.013 48.496 43.213 ;
 RECT 48.272 43.013 48.328 43.213 ;
 RECT 47.768 43.147 47.824 43.347 ;
 RECT 47.768 40.627 47.824 40.827 ;
 RECT 49.532 40.703 49.588 40.903 ;
 RECT 47.768 41.887 47.824 42.087 ;
 RECT 47.6 41.199 47.656 41.399 ;
 RECT 49.28 41.4035 49.336 41.6035 ;
 RECT 46.928 41.188 46.984 41.388 ;
 RECT 47.432 41.137 47.488 41.337 ;
 RECT 47.264 41.188 47.32 41.388 ;
 RECT 46.592 41.218 46.648 41.418 ;
 RECT 46.76 41.218 46.816 41.418 ;
 RECT 47.096 41.188 47.152 41.388 ;
 END
 END vss.gds3571
 PIN vss.gds3572
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.542 43.8995 51.598 44.0995 ;
 END
 END vss.gds3572
 PIN vss.gds3573
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 41.796 50.918 41.996 ;
 END
 END vss.gds3573
 PIN vss.gds3574
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.638 41.3235 52.698 41.5235 ;
 END
 END vss.gds3574
 PIN vss.gds3575
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.806 41.3235 52.866 41.5235 ;
 END
 END vss.gds3575
 PIN vss.gds3576
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.142 41.3235 53.202 41.5235 ;
 END
 END vss.gds3576
 PIN vss.gds3577
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.31 41.3235 53.37 41.5235 ;
 END
 END vss.gds3577
 PIN vss.gds3578
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.478 41.3235 53.538 41.5235 ;
 END
 END vss.gds3578
 PIN vss.gds3579
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.814 41.3235 53.874 41.5235 ;
 END
 END vss.gds3579
 PIN vss.gds3580
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.982 41.3235 54.042 41.5235 ;
 END
 END vss.gds3580
 PIN vss.gds3581
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.15 41.3235 54.21 41.5235 ;
 END
 END vss.gds3581
 PIN vss.gds3582
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.486 41.3235 54.546 41.5235 ;
 END
 END vss.gds3582
 PIN vss.gds3583
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.654 41.3235 54.714 41.5235 ;
 END
 END vss.gds3583
 PIN vss.gds3584
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.822 41.3235 54.882 41.5235 ;
 END
 END vss.gds3584
 PIN vss.gds3585
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 42.9595 55.05 43.1595 ;
 END
 END vss.gds3585
 PIN vss.gds3586
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.158 41.3235 55.218 41.5235 ;
 END
 END vss.gds3586
 PIN vss.gds3587
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 42.9595 54.378 43.1595 ;
 END
 END vss.gds3587
 PIN vss.gds3588
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 42.9595 53.706 43.1595 ;
 END
 END vss.gds3588
 PIN vss.gds3589
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.47 41.3235 52.53 41.5235 ;
 END
 END vss.gds3589
 PIN vss.gds3590
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 44.7555 51.418 44.9555 ;
 END
 END vss.gds3590
 PIN vss.gds3591
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.09 41.107 52.13 41.307 ;
 END
 END vss.gds3591
 PIN vss.gds3592
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 43.0465 51.098 43.2465 ;
 END
 END vss.gds3592
 PIN vss.gds3593
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 42.9595 53.034 43.1595 ;
 END
 END vss.gds3593
 PIN vss.gds3594
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 43.1235 51.938 43.3235 ;
 END
 END vss.gds3594
 PIN vss.gds3595
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 43.2305 50.594 43.4305 ;
 END
 END vss.gds3595
 PIN vss.gds3596
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 42.925 52.362 43.125 ;
 END
 END vss.gds3596
 PIN vss.gds3597
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 50.624 44.96 50.68 45.113 ;
 RECT 50.624 43.7 50.68 43.853 ;
 RECT 50.624 41.18 50.68 41.333 ;
 RECT 50.624 42.44 50.68 42.593 ;
 RECT 50.456 44.5835 50.512 44.7835 ;
 RECT 50.96 44.3315 51.016 44.5315 ;
 RECT 50.456 40.8035 50.512 41.0035 ;
 RECT 50.96 40.5515 51.016 40.7515 ;
 RECT 50.96 43.0715 51.016 43.2715 ;
 RECT 50.456 43.3235 50.512 43.5235 ;
 RECT 50.456 42.0635 50.512 42.2635 ;
 RECT 50.96 41.8115 51.016 42.0115 ;
 RECT 51.968 41.218 52.024 41.418 ;
 RECT 51.8 41.2255 51.856 41.4255 ;
 RECT 51.632 41.218 51.688 41.418 ;
 RECT 51.464 41.218 51.52 41.418 ;
 RECT 51.296 41.218 51.352 41.418 ;
 RECT 51.128 41.333 51.184 41.533 ;
 RECT 52.136 41.218 52.192 41.418 ;
 END
 END vss.gds3597
 PIN vss.gds3598
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 42.9595 60.174 43.1595 ;
 END
 END vss.gds3598
 PIN vss.gds3599
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.946 41.3235 60.006 41.5235 ;
 END
 END vss.gds3599
 PIN vss.gds3600
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.778 41.3235 59.838 41.5235 ;
 END
 END vss.gds3600
 PIN vss.gds3601
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.61 41.3235 59.67 41.5235 ;
 END
 END vss.gds3601
 PIN vss.gds3602
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 42.9595 59.502 43.1595 ;
 END
 END vss.gds3602
 PIN vss.gds3603
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.274 41.3235 59.334 41.5235 ;
 END
 END vss.gds3603
 PIN vss.gds3604
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.106 41.3235 59.166 41.5235 ;
 END
 END vss.gds3604
 PIN vss.gds3605
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.938 41.3235 58.998 41.5235 ;
 END
 END vss.gds3605
 PIN vss.gds3606
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 42.9595 58.83 43.1595 ;
 END
 END vss.gds3606
 PIN vss.gds3607
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.602 41.3235 58.662 41.5235 ;
 END
 END vss.gds3607
 PIN vss.gds3608
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.434 41.3235 58.494 41.5235 ;
 END
 END vss.gds3608
 PIN vss.gds3609
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.266 41.3235 58.326 41.5235 ;
 END
 END vss.gds3609
 PIN vss.gds3610
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.326 41.3235 55.386 41.5235 ;
 END
 END vss.gds3610
 PIN vss.gds3611
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.494 41.3235 55.554 41.5235 ;
 END
 END vss.gds3611
 PIN vss.gds3612
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.83 41.3235 55.89 41.5235 ;
 END
 END vss.gds3612
 PIN vss.gds3613
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.998 41.3235 56.058 41.5235 ;
 END
 END vss.gds3613
 PIN vss.gds3614
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.166 41.3235 56.226 41.5235 ;
 END
 END vss.gds3614
 PIN vss.gds3615
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.502 41.3235 56.562 41.5235 ;
 END
 END vss.gds3615
 PIN vss.gds3616
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.67 41.3235 56.73 41.5235 ;
 END
 END vss.gds3616
 PIN vss.gds3617
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.838 41.3235 56.898 41.5235 ;
 END
 END vss.gds3617
 PIN vss.gds3618
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.342 41.3235 57.402 41.5235 ;
 END
 END vss.gds3618
 PIN vss.gds3619
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.51 41.3235 57.57 41.5235 ;
 END
 END vss.gds3619
 PIN vss.gds3620
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 42.9595 55.722 43.1595 ;
 END
 END vss.gds3620
 PIN vss.gds3621
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 42.9595 56.394 43.1595 ;
 END
 END vss.gds3621
 PIN vss.gds3622
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.174 41.3235 57.234 41.5235 ;
 END
 END vss.gds3622
 PIN vss.gds3623
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 42.9595 57.738 43.1595 ;
 END
 END vss.gds3623
 PIN vss.gds3624
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 42.9595 57.066 43.1595 ;
 END
 END vss.gds3624
 PIN vss.gds3625
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 58.016 44.42 58.072 44.62 ;
 RECT 58.016 41.9 58.072 42.1 ;
 RECT 58.016 40.64 58.072 40.84 ;
 RECT 58.016 43.16 58.072 43.36 ;
 RECT 57.848 43.09 57.904 43.29 ;
 END
 END vss.gds3625
 PIN vss.gds3626
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 40.982 65.054 41.182 ;
 END
 END vss.gds3626
 PIN vss.gds3627
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 42.242 65.054 42.442 ;
 END
 END vss.gds3627
 PIN vss.gds3628
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 43.502 65.054 43.702 ;
 END
 END vss.gds3628
 PIN vss.gds3629
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 42.0095 64.214 42.2095 ;
 END
 END vss.gds3629
 PIN vss.gds3630
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.418 44.316 64.474 44.516 ;
 END
 END vss.gds3630
 PIN vss.gds3631
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 42.925 63.534 43.125 ;
 END
 END vss.gds3631
 PIN vss.gds3632
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.306 41.3235 63.366 41.5235 ;
 END
 END vss.gds3632
 PIN vss.gds3633
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.138 41.3235 63.198 41.5235 ;
 END
 END vss.gds3633
 PIN vss.gds3634
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.97 41.3235 63.03 41.5235 ;
 END
 END vss.gds3634
 PIN vss.gds3635
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 42.9595 62.862 43.1595 ;
 END
 END vss.gds3635
 PIN vss.gds3636
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.634 41.3235 62.694 41.5235 ;
 END
 END vss.gds3636
 PIN vss.gds3637
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.466 41.3235 62.526 41.5235 ;
 END
 END vss.gds3637
 PIN vss.gds3638
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.298 41.3235 62.358 41.5235 ;
 END
 END vss.gds3638
 PIN vss.gds3639
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 42.9595 62.19 43.1595 ;
 END
 END vss.gds3639
 PIN vss.gds3640
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.962 41.3235 62.022 41.5235 ;
 END
 END vss.gds3640
 PIN vss.gds3641
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.794 41.3235 61.854 41.5235 ;
 END
 END vss.gds3641
 PIN vss.gds3642
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.626 41.3235 61.686 41.5235 ;
 END
 END vss.gds3642
 PIN vss.gds3643
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 42.9595 61.518 43.1595 ;
 END
 END vss.gds3643
 PIN vss.gds3644
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.29 41.3235 61.35 41.5235 ;
 END
 END vss.gds3644
 PIN vss.gds3645
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.122 41.3235 61.182 41.5235 ;
 END
 END vss.gds3645
 PIN vss.gds3646
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.954 41.3235 61.014 41.5235 ;
 END
 END vss.gds3646
 PIN vss.gds3647
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 42.9595 60.846 43.1595 ;
 END
 END vss.gds3647
 PIN vss.gds3648
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.618 41.3235 60.678 41.5235 ;
 END
 END vss.gds3648
 PIN vss.gds3649
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.45 41.3235 60.51 41.5235 ;
 END
 END vss.gds3649
 PIN vss.gds3650
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.282 41.3235 60.342 41.5235 ;
 END
 END vss.gds3650
 PIN vss.gds3651
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 43.1235 63.974 43.3235 ;
 END
 END vss.gds3651
 PIN vss.gds3652
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 43.627 63.746 43.827 ;
 END
 END vss.gds3652
 PIN vss.gds3653
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 44.762 65.054 44.962 ;
 END
 END vss.gds3653
 PIN vss.gds3654
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 42.9595 64.814 43.1595 ;
 END
 END vss.gds3654
 PIN vss.gds3655
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 65.156 44.94 65.212 45.113 ;
 RECT 65.156 43.68 65.212 43.853 ;
 RECT 65.156 41.16 65.212 41.333 ;
 RECT 65.156 42.42 65.212 42.593 ;
 RECT 64.82 44.407 64.876 44.607 ;
 RECT 64.82 43.147 64.876 43.347 ;
 RECT 64.82 41.887 64.876 42.087 ;
 RECT 64.82 40.627 64.876 40.827 ;
 RECT 64.652 41.199 64.708 41.399 ;
 RECT 63.98 41.188 64.036 41.388 ;
 RECT 63.812 41.218 63.868 41.418 ;
 RECT 64.484 41.137 64.54 41.337 ;
 RECT 64.316 41.188 64.372 41.388 ;
 RECT 63.644 41.218 63.7 41.418 ;
 RECT 64.148 41.188 64.204 41.388 ;
 END
 END vss.gds3655
 PIN vss.gds3656
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 42.282 66.026 42.482 ;
 END
 END vss.gds3656
 PIN vss.gds3657
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 41.022 66.026 41.222 ;
 END
 END vss.gds3657
 PIN vss.gds3658
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 43.542 66.026 43.742 ;
 END
 END vss.gds3658
 PIN vss.gds3659
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 44.802 66.026 45.002 ;
 END
 END vss.gds3659
 PIN vss.gds3660
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 45 66.574 45.2 ;
 END
 END vss.gds3660
 PIN vss.gds3661
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.594 43.8995 68.65 44.0995 ;
 END
 END vss.gds3661
 PIN vss.gds3662
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 43.0465 68.15 43.2465 ;
 END
 END vss.gds3662
 PIN vss.gds3663
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.858 41.3235 69.918 41.5235 ;
 END
 END vss.gds3663
 PIN vss.gds3664
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.194 41.3235 70.254 41.5235 ;
 END
 END vss.gds3664
 PIN vss.gds3665
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.142 41.107 69.182 41.307 ;
 END
 END vss.gds3665
 PIN vss.gds3666
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 44.257 67.302 44.457 ;
 END
 END vss.gds3666
 PIN vss.gds3667
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 42.997 67.302 43.197 ;
 END
 END vss.gds3667
 PIN vss.gds3668
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 41.737 67.302 41.937 ;
 END
 END vss.gds3668
 PIN vss.gds3669
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 40.477 67.302 40.677 ;
 END
 END vss.gds3669
 PIN vss.gds3670
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 41.796 67.97 41.996 ;
 END
 END vss.gds3670
 PIN vss.gds3671
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.69 41.3235 69.75 41.5235 ;
 END
 END vss.gds3671
 PIN vss.gds3672
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 43.128 66.318 43.328 ;
 END
 END vss.gds3672
 PIN vss.gds3673
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.522 41.3235 69.582 41.5235 ;
 END
 END vss.gds3673
 PIN vss.gds3674
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 44.7555 68.47 44.9555 ;
 END
 END vss.gds3674
 PIN vss.gds3675
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 42.9595 70.086 43.1595 ;
 END
 END vss.gds3675
 PIN vss.gds3676
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 43.128 66.998 43.328 ;
 END
 END vss.gds3676
 PIN vss.gds3677
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 43.128 65.654 43.328 ;
 END
 END vss.gds3677
 PIN vss.gds3678
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 43.2305 67.646 43.4305 ;
 END
 END vss.gds3678
 PIN vss.gds3679
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 43.1235 68.99 43.3235 ;
 END
 END vss.gds3679
 PIN vss.gds3680
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 42.925 69.414 43.125 ;
 END
 END vss.gds3680
 PIN vss.gds3681
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 67.676 44.96 67.732 45.113 ;
 RECT 65.324 44.913 65.38 45.113 ;
 RECT 66.92 44.957 66.976 45.122 ;
 RECT 66.752 44.957 66.808 45.122 ;
 RECT 65.996 44.957 66.052 45.122 ;
 RECT 65.828 44.957 65.884 45.122 ;
 RECT 67.676 43.7 67.732 43.853 ;
 RECT 65.324 43.653 65.38 43.853 ;
 RECT 66.92 43.697 66.976 43.862 ;
 RECT 66.752 43.697 66.808 43.862 ;
 RECT 65.996 43.697 66.052 43.862 ;
 RECT 65.828 43.697 65.884 43.862 ;
 RECT 67.676 41.18 67.732 41.333 ;
 RECT 65.324 41.133 65.38 41.333 ;
 RECT 66.92 41.177 66.976 41.342 ;
 RECT 66.752 41.177 66.808 41.342 ;
 RECT 65.996 41.177 66.052 41.342 ;
 RECT 65.828 41.177 65.884 41.342 ;
 RECT 67.676 42.44 67.732 42.593 ;
 RECT 65.324 42.393 65.38 42.593 ;
 RECT 66.92 42.437 66.976 42.602 ;
 RECT 66.752 42.437 66.808 42.602 ;
 RECT 65.996 42.437 66.052 42.602 ;
 RECT 65.828 42.437 65.884 42.602 ;
 RECT 66.752 41.404 66.808 41.604 ;
 RECT 67.004 41.407 67.06 41.607 ;
 RECT 66.752 42.664 66.808 42.864 ;
 RECT 67.004 42.667 67.06 42.867 ;
 RECT 66.752 43.924 66.808 44.124 ;
 RECT 67.004 43.927 67.06 44.127 ;
 RECT 66.752 45.184 66.808 45.384 ;
 RECT 67.004 45.187 67.06 45.387 ;
 RECT 65.492 44.273 65.548 44.473 ;
 RECT 65.324 44.273 65.38 44.473 ;
 RECT 66.164 44.483 66.22 44.683 ;
 RECT 66.584 44.483 66.64 44.683 ;
 RECT 67.508 44.5835 67.564 44.7835 ;
 RECT 68.012 44.3315 68.068 44.5315 ;
 RECT 66.164 41.963 66.22 42.163 ;
 RECT 65.492 41.753 65.548 41.953 ;
 RECT 65.324 41.753 65.38 41.953 ;
 RECT 67.508 42.0635 67.564 42.2635 ;
 RECT 68.012 41.8115 68.068 42.0115 ;
 RECT 68.012 43.0715 68.068 43.2715 ;
 RECT 67.508 43.3235 67.564 43.5235 ;
 RECT 66.164 43.223 66.22 43.423 ;
 RECT 66.584 43.223 66.64 43.423 ;
 RECT 65.492 43.013 65.548 43.213 ;
 RECT 65.324 43.013 65.38 43.213 ;
 RECT 66.584 41.963 66.64 42.163 ;
 RECT 68.012 40.5515 68.068 40.7515 ;
 RECT 67.508 40.8035 67.564 41.0035 ;
 RECT 66.164 40.703 66.22 40.903 ;
 RECT 66.584 40.703 66.64 40.903 ;
 RECT 65.492 40.493 65.548 40.693 ;
 RECT 65.324 40.493 65.38 40.693 ;
 RECT 66.332 41.4035 66.388 41.6035 ;
 RECT 69.02 41.218 69.076 41.418 ;
 RECT 68.852 41.2255 68.908 41.4255 ;
 RECT 68.684 41.218 68.74 41.418 ;
 RECT 68.516 41.218 68.572 41.418 ;
 RECT 68.348 41.218 68.404 41.418 ;
 RECT 69.188 41.218 69.244 41.418 ;
 RECT 68.18 41.333 68.236 41.533 ;
 END
 END vss.gds3681
 PIN vss.gds3682
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.362 41.3235 70.422 41.5235 ;
 END
 END vss.gds3682
 PIN vss.gds3683
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.53 41.3235 70.59 41.5235 ;
 END
 END vss.gds3683
 PIN vss.gds3684
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.866 41.3235 70.926 41.5235 ;
 END
 END vss.gds3684
 PIN vss.gds3685
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.034 41.3235 71.094 41.5235 ;
 END
 END vss.gds3685
 PIN vss.gds3686
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.202 41.3235 71.262 41.5235 ;
 END
 END vss.gds3686
 PIN vss.gds3687
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 42.9595 71.43 43.1595 ;
 END
 END vss.gds3687
 PIN vss.gds3688
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.538 41.3235 71.598 41.5235 ;
 END
 END vss.gds3688
 PIN vss.gds3689
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.706 41.3235 71.766 41.5235 ;
 END
 END vss.gds3689
 PIN vss.gds3690
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.874 41.3235 71.934 41.5235 ;
 END
 END vss.gds3690
 PIN vss.gds3691
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 42.9595 72.102 43.1595 ;
 END
 END vss.gds3691
 PIN vss.gds3692
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.21 41.3235 72.27 41.5235 ;
 END
 END vss.gds3692
 PIN vss.gds3693
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.378 41.3235 72.438 41.5235 ;
 END
 END vss.gds3693
 PIN vss.gds3694
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.546 41.3235 72.606 41.5235 ;
 END
 END vss.gds3694
 PIN vss.gds3695
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 42.9595 72.774 43.1595 ;
 END
 END vss.gds3695
 PIN vss.gds3696
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.882 41.3235 72.942 41.5235 ;
 END
 END vss.gds3696
 PIN vss.gds3697
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.05 41.3235 73.11 41.5235 ;
 END
 END vss.gds3697
 PIN vss.gds3698
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.554 41.3235 73.614 41.5235 ;
 END
 END vss.gds3698
 PIN vss.gds3699
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.722 41.3235 73.782 41.5235 ;
 END
 END vss.gds3699
 PIN vss.gds3700
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.89 41.3235 73.95 41.5235 ;
 END
 END vss.gds3700
 PIN vss.gds3701
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.394 41.3235 74.454 41.5235 ;
 END
 END vss.gds3701
 PIN vss.gds3702
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.218 41.3235 73.278 41.5235 ;
 END
 END vss.gds3702
 PIN vss.gds3703
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.562 41.3235 74.622 41.5235 ;
 END
 END vss.gds3703
 PIN vss.gds3704
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.226 41.3235 74.286 41.5235 ;
 END
 END vss.gds3704
 PIN vss.gds3705
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 42.9595 70.758 43.1595 ;
 END
 END vss.gds3705
 PIN vss.gds3706
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 42.9595 73.446 43.1595 ;
 END
 END vss.gds3706
 PIN vss.gds3707
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 42.9595 74.118 43.1595 ;
 END
 END vss.gds3707
 PIN vss.gds3708
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 42.9595 74.79 43.1595 ;
 END
 END vss.gds3708
 PIN vss.gds3709
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 45.517 2.962 45.717 ;
 END
 END vss.gds3709
 PIN vss.gds3710
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 48.037 2.962 48.237 ;
 END
 END vss.gds3710
 PIN vss.gds3711
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.906 46.777 2.962 46.977 ;
 END
 END vss.gds3711
 PIN vss.gds3712
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 48.726 3.142 48.926 ;
 END
 END vss.gds3712
 PIN vss.gds3713
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 46.376 3.142 46.576 ;
 END
 END vss.gds3713
 PIN vss.gds3714
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.442 45.741 4.482 45.941 ;
 END
 END vss.gds3714
 PIN vss.gds3715
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.286 46.147 3.326 46.347 ;
 END
 END vss.gds3715
 PIN vss.gds3716
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.754 47.407 3.794 47.607 ;
 END
 END vss.gds3716
 PIN vss.gds3717
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.57 45.944 4.61 46.144 ;
 END
 END vss.gds3717
 PIN vss.gds3718
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.414 46.423 3.454 46.623 ;
 END
 END vss.gds3718
 PIN vss.gds3719
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.842 45.741 4.882 45.941 ;
 END
 END vss.gds3719
 PIN vss.gds3720
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.034 47.407 5.074 47.607 ;
 END
 END vss.gds3720
 PIN vss.gds3721
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.562 46.423 3.602 46.623 ;
 END
 END vss.gds3721
 PIN vss.gds3722
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.066 47.636 3.142 47.836 ;
 END
 END vss.gds3722
 PIN vss.gds3723
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.882 47.001 0.942 47.201 ;
 END
 END vss.gds3723
 PIN vss.gds3724
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 4.154 47.407 4.194 47.607 ;
 END
 END vss.gds3724
 PIN vss.gds3725
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.678 47.1015 0.718 47.3015 ;
 END
 END vss.gds3725
 PIN vss.gds3726
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.572 47.202 0.602 47.402 ;
 END
 END vss.gds3726
 PIN vss.gds3727
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.066 47.1965 2.122 47.3965 ;
 END
 END vss.gds3727
 PIN vss.gds3728
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.242 47.545 1.282 47.745 ;
 END
 END vss.gds3728
 PIN vss.gds3729
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 1.386 47.448 1.462 47.648 ;
 END
 END vss.gds3729
 PIN vss.gds3730
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 2.226 47.032 2.302 47.232 ;
 END
 END vss.gds3730
 PIN vss.gds3731
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 3.946 47.3035 4.002 47.5035 ;
 END
 END vss.gds3731
 PIN vss.gds3732
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.226 47.3035 5.282 47.5035 ;
 END
 END vss.gds3732
 PIN vss.gds3733
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 0.234 47.78 0.29 47.98 ;
 END
 END vss.gds3733
 PIN vss.gds3734
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 2.576 45.5175 2.632 45.7175 ;
 RECT 2.408 45.5175 2.464 45.7175 ;
 RECT 2.996 45.5175 3.052 45.7175 ;
 RECT 3.332 45.609 3.388 45.809 ;
 RECT 2.408 46.7775 2.464 46.9775 ;
 RECT 2.576 46.7775 2.632 46.9775 ;
 RECT 2.996 46.7775 3.052 46.9775 ;
 RECT 3.332 46.869 3.388 47.069 ;
 RECT 3.5 46.8255 3.556 47.0255 ;
 RECT 0.98 46.6925 1.036 46.8925 ;
 RECT 2.072 46.693 2.128 46.893 ;
 RECT 2.576 48.0375 2.632 48.2375 ;
 RECT 2.408 48.0375 2.464 48.2375 ;
 RECT 2.996 48.0375 3.052 48.2375 ;
 RECT 3.332 48.129 3.388 48.329 ;
 RECT 0.812 45.609 0.868 45.809 ;
 RECT 3.5 48.0855 3.556 48.2855 ;
 RECT 0.98 47.9525 1.036 48.1525 ;
 RECT 2.072 47.953 2.128 48.153 ;
 RECT 0.392 48.043 0.448 48.243 ;
 RECT 0.812 48.129 0.868 48.329 ;
 RECT 0.644 48.043 0.7 48.243 ;
 RECT 1.232 48.043 1.288 48.243 ;
 RECT 1.4 48.043 1.456 48.243 ;
 RECT 1.568 48.043 1.624 48.243 ;
 RECT 1.82 48.043 1.876 48.243 ;
 RECT 2.24 48.043 2.296 48.243 ;
 RECT 2.744 47.953 2.8 48.153 ;
 RECT 3.164 48.043 3.22 48.243 ;
 RECT 3.5 45.5655 3.556 45.7655 ;
 RECT 0.392 45.523 0.448 45.723 ;
 RECT 0.644 45.523 0.7 45.723 ;
 RECT 1.232 45.523 1.288 45.723 ;
 RECT 1.4 45.523 1.456 45.723 ;
 RECT 1.568 45.523 1.624 45.723 ;
 RECT 1.82 45.523 1.876 45.723 ;
 RECT 3.164 45.523 3.22 45.723 ;
 RECT 2.24 45.523 2.296 45.723 ;
 RECT 3.92 48.043 3.976 48.243 ;
 RECT 3.752 48.313 3.808 48.513 ;
 RECT 4.508 48.2425 4.564 48.4425 ;
 RECT 0.392 46.783 0.448 46.983 ;
 RECT 0.812 46.869 0.868 47.069 ;
 RECT 0.644 46.783 0.7 46.983 ;
 RECT 1.232 46.783 1.288 46.983 ;
 RECT 1.4 46.783 1.456 46.983 ;
 RECT 1.568 46.783 1.624 46.983 ;
 RECT 1.82 46.783 1.876 46.983 ;
 RECT 2.24 46.783 2.296 46.983 ;
 RECT 2.744 46.693 2.8 46.893 ;
 RECT 3.164 46.783 3.22 46.983 ;
 RECT 3.92 46.783 3.976 46.983 ;
 RECT 3.752 47.053 3.808 47.253 ;
 RECT 4.508 46.9825 4.564 47.1825 ;
 RECT 3.92 45.523 3.976 45.723 ;
 RECT 3.752 45.793 3.808 45.993 ;
 RECT 4.508 45.7225 4.564 45.9225 ;
 END
 END vss.gds3734
 PIN vss.gds3735
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.134 46.3635 10.194 46.5635 ;
 END
 END vss.gds3735
 PIN vss.gds3736
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.966 46.3635 10.026 46.5635 ;
 END
 END vss.gds3736
 PIN vss.gds3737
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.798 46.3635 9.858 46.5635 ;
 END
 END vss.gds3737
 PIN vss.gds3738
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.462 46.3635 9.522 46.5635 ;
 END
 END vss.gds3738
 PIN vss.gds3739
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.294 46.3635 9.354 46.5635 ;
 END
 END vss.gds3739
 PIN vss.gds3740
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.79 46.3635 8.85 46.5635 ;
 END
 END vss.gds3740
 PIN vss.gds3741
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.622 46.3635 8.682 46.5635 ;
 END
 END vss.gds3741
 PIN vss.gds3742
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.454 46.3635 8.514 46.5635 ;
 END
 END vss.gds3742
 PIN vss.gds3743
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.118 46.3635 8.178 46.5635 ;
 END
 END vss.gds3743
 PIN vss.gds3744
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.95 46.3635 8.01 46.5635 ;
 END
 END vss.gds3744
 PIN vss.gds3745
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.782 46.3635 7.842 46.5635 ;
 END
 END vss.gds3745
 PIN vss.gds3746
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.126 46.3635 9.186 46.5635 ;
 END
 END vss.gds3746
 PIN vss.gds3747
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.446 46.3635 7.506 46.5635 ;
 END
 END vss.gds3747
 PIN vss.gds3748
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.278 46.3635 7.338 46.5635 ;
 END
 END vss.gds3748
 PIN vss.gds3749
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 9.63 47.128 9.69 47.328 ;
 END
 END vss.gds3749
 PIN vss.gds3750
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.958 47.128 9.018 47.328 ;
 END
 END vss.gds3750
 PIN vss.gds3751
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.11 46.3635 7.17 46.5635 ;
 END
 END vss.gds3751
 PIN vss.gds3752
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.138 47.204 6.178 47.404 ;
 END
 END vss.gds3752
 PIN vss.gds3753
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.434 47.407 5.474 47.607 ;
 END
 END vss.gds3753
 PIN vss.gds3754
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 8.286 47.128 8.346 47.328 ;
 END
 END vss.gds3754
 PIN vss.gds3755
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 7.614 47.128 7.674 47.328 ;
 END
 END vss.gds3755
 PIN vss.gds3756
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.69 47.407 5.73 47.607 ;
 END
 END vss.gds3756
 PIN vss.gds3757
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 5.946 47.407 5.986 47.607 ;
 END
 END vss.gds3757
 PIN vss.gds3758
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 6.394 46.962 6.434 47.162 ;
 END
 END vss.gds3758
 PIN vss.gds3759
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 6.692 48.186 6.748 48.386 ;
 RECT 6.524 48.036 6.58 48.236 ;
 RECT 6.608 48.313 6.664 48.513 ;
 RECT 6.608 47.053 6.664 47.253 ;
 RECT 6.524 46.776 6.58 46.976 ;
 RECT 6.692 46.926 6.748 47.126 ;
 RECT 6.692 45.666 6.748 45.866 ;
 RECT 6.524 45.516 6.58 45.716 ;
 RECT 6.608 45.793 6.664 45.993 ;
 END
 END vss.gds3759
 PIN vss.gds3760
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 47.322 14.87 47.522 ;
 END
 END vss.gds3760
 PIN vss.gds3761
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 48.542 13.898 48.742 ;
 END
 END vss.gds3761
 PIN vss.gds3762
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 48.582 14.87 48.782 ;
 END
 END vss.gds3762
 PIN vss.gds3763
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 46.022 13.898 46.222 ;
 END
 END vss.gds3763
 PIN vss.gds3764
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.83 46.062 14.87 46.262 ;
 END
 END vss.gds3764
 PIN vss.gds3765
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.15 46.3635 12.21 46.5635 ;
 END
 END vss.gds3765
 PIN vss.gds3766
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.982 46.3635 12.042 46.5635 ;
 END
 END vss.gds3766
 PIN vss.gds3767
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.814 46.3635 11.874 46.5635 ;
 END
 END vss.gds3767
 PIN vss.gds3768
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.478 46.3635 11.538 46.5635 ;
 END
 END vss.gds3768
 PIN vss.gds3769
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.31 46.3635 11.37 46.5635 ;
 END
 END vss.gds3769
 PIN vss.gds3770
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.142 46.3635 11.202 46.5635 ;
 END
 END vss.gds3770
 PIN vss.gds3771
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.806 46.3635 10.866 46.5635 ;
 END
 END vss.gds3771
 PIN vss.gds3772
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.638 46.3635 10.698 46.5635 ;
 END
 END vss.gds3772
 PIN vss.gds3773
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.47 46.3635 10.53 46.5635 ;
 END
 END vss.gds3773
 PIN vss.gds3774
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.002 46.728 13.058 46.928 ;
 END
 END vss.gds3774
 PIN vss.gds3775
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.262 47.937 13.318 48.137 ;
 END
 END vss.gds3775
 PIN vss.gds3776
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 11.646 47.128 11.706 47.328 ;
 END
 END vss.gds3776
 PIN vss.gds3777
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.974 47.128 11.034 47.328 ;
 END
 END vss.gds3777
 PIN vss.gds3778
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 10.302 47.128 10.362 47.328 ;
 END
 END vss.gds3778
 PIN vss.gds3779
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.102 47.283 15.162 47.483 ;
 END
 END vss.gds3779
 PIN vss.gds3780
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.842 47.282 13.898 47.482 ;
 END
 END vss.gds3780
 PIN vss.gds3781
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 14.422 47.283 14.498 47.483 ;
 END
 END vss.gds3781
 PIN vss.gds3782
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 13.582 47.128 13.658 47.328 ;
 END
 END vss.gds3782
 PIN vss.gds3783
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.318 47.1405 12.378 47.3405 ;
 END
 END vss.gds3783
 PIN vss.gds3784
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.55 47.407 12.59 47.607 ;
 END
 END vss.gds3784
 PIN vss.gds3785
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 12.742 47.157 12.818 47.357 ;
 END
 END vss.gds3785
 PIN vss.gds3786
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 14 48.72 14.056 48.893 ;
 RECT 14.168 48.693 14.224 48.893 ;
 RECT 14 47.46 14.056 47.633 ;
 RECT 14.168 47.433 14.224 47.633 ;
 RECT 14 46.2 14.056 46.373 ;
 RECT 14.168 46.173 14.224 46.373 ;
 RECT 14.336 45.533 14.392 45.733 ;
 RECT 14.168 45.533 14.224 45.733 ;
 RECT 15.008 45.743 15.064 45.943 ;
 RECT 14.84 46.217 14.896 46.382 ;
 RECT 14.672 46.217 14.728 46.382 ;
 RECT 13.664 45.667 13.72 45.867 ;
 RECT 14.336 46.793 14.392 46.993 ;
 RECT 14.168 46.793 14.224 46.993 ;
 RECT 13.664 46.927 13.72 47.127 ;
 RECT 14.84 47.477 14.896 47.642 ;
 RECT 14.672 47.477 14.728 47.642 ;
 RECT 15.008 47.003 15.064 47.203 ;
 RECT 15.008 48.263 15.064 48.463 ;
 RECT 14.84 48.737 14.896 48.902 ;
 RECT 14.672 48.737 14.728 48.902 ;
 RECT 14.336 48.053 14.392 48.253 ;
 RECT 14.168 48.053 14.224 48.253 ;
 RECT 13.664 48.187 13.72 48.387 ;
 RECT 15.176 48.83 15.232 49.03 ;
 RECT 15.176 46.3665 15.232 46.5665 ;
 RECT 12.824 48.767 12.88 48.967 ;
 RECT 12.824 46.1645 12.88 46.3645 ;
 RECT 13.496 46.239 13.552 46.439 ;
 RECT 13.328 48.767 13.384 48.967 ;
 RECT 13.328 46.1045 13.384 46.3045 ;
 RECT 13.16 48.767 13.216 48.967 ;
 RECT 13.16 46.1645 13.216 46.3645 ;
 RECT 12.488 48.767 12.544 48.967 ;
 RECT 12.488 46.2015 12.544 46.4015 ;
 RECT 12.992 48.767 13.048 48.967 ;
 RECT 12.992 46.1645 13.048 46.3645 ;
 RECT 12.656 48.767 12.712 48.967 ;
 RECT 12.656 46.2015 12.712 46.4015 ;
 END
 END vss.gds3786
 PIN vss.gds3787
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.378 48.15 15.418 48.35 ;
 END
 END vss.gds3787
 PIN vss.gds3788
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.438 47.6795 17.494 47.8795 ;
 END
 END vss.gds3788
 PIN vss.gds3789
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 48.037 16.146 48.237 ;
 END
 END vss.gds3789
 PIN vss.gds3790
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 46.777 16.146 46.977 ;
 END
 END vss.gds3790
 PIN vss.gds3791
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.214 47.128 20.274 47.328 ;
 END
 END vss.gds3791
 PIN vss.gds3792
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.1 45.517 16.146 45.717 ;
 END
 END vss.gds3792
 PIN vss.gds3793
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.702 46.3635 18.762 46.5635 ;
 END
 END vss.gds3793
 PIN vss.gds3794
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.038 46.3635 19.098 46.5635 ;
 END
 END vss.gds3794
 PIN vss.gds3795
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.206 46.3635 19.266 46.5635 ;
 END
 END vss.gds3795
 PIN vss.gds3796
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.374 46.3635 19.434 46.5635 ;
 END
 END vss.gds3796
 PIN vss.gds3797
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.71 46.3635 19.77 46.5635 ;
 END
 END vss.gds3797
 PIN vss.gds3798
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.878 46.3635 19.938 46.5635 ;
 END
 END vss.gds3798
 PIN vss.gds3799
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.534 46.3635 18.594 46.5635 ;
 END
 END vss.gds3799
 PIN vss.gds3800
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.758 46.6495 16.814 46.8495 ;
 END
 END vss.gds3800
 PIN vss.gds3801
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.366 46.3635 18.426 46.5635 ;
 END
 END vss.gds3801
 PIN vss.gds3802
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.258 48.039 17.314 48.239 ;
 END
 END vss.gds3802
 PIN vss.gds3803
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.986 46.147 18.026 46.347 ;
 END
 END vss.gds3803
 PIN vss.gds3804
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.87 47.128 18.93 47.328 ;
 END
 END vss.gds3804
 PIN vss.gds3805
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 19.542 47.128 19.602 47.328 ;
 END
 END vss.gds3805
 PIN vss.gds3806
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.918 47.2205 16.994 47.4205 ;
 END
 END vss.gds3806
 PIN vss.gds3807
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.046 46.3635 20.106 46.5635 ;
 END
 END vss.gds3807
 PIN vss.gds3808
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 15.766 47.283 15.842 47.483 ;
 END
 END vss.gds3808
 PIN vss.gds3809
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 18.198 47.1405 18.258 47.3405 ;
 END
 END vss.gds3809
 PIN vss.gds3810
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 17.758 47.157 17.834 47.357 ;
 END
 END vss.gds3810
 PIN vss.gds3811
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 16.414 47.1965 16.49 47.3965 ;
 END
 END vss.gds3811
 PIN vss.gds3812
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 15.596 47.704 15.652 47.904 ;
 RECT 15.848 47.707 15.904 47.907 ;
 RECT 16.52 48.74 16.576 48.893 ;
 RECT 15.764 48.737 15.82 48.902 ;
 RECT 15.596 48.737 15.652 48.902 ;
 RECT 15.596 46.444 15.652 46.644 ;
 RECT 15.848 46.447 15.904 46.647 ;
 RECT 16.52 47.48 16.576 47.633 ;
 RECT 16.52 46.22 16.576 46.373 ;
 RECT 15.764 46.217 15.82 46.382 ;
 RECT 15.596 46.217 15.652 46.382 ;
 RECT 15.428 45.743 15.484 45.943 ;
 RECT 16.352 45.8435 16.408 46.0435 ;
 RECT 16.856 45.5915 16.912 45.7915 ;
 RECT 16.352 47.1035 16.408 47.3035 ;
 RECT 16.856 46.8515 16.912 47.0515 ;
 RECT 15.764 47.477 15.82 47.642 ;
 RECT 15.596 47.477 15.652 47.642 ;
 RECT 15.428 47.003 15.484 47.203 ;
 RECT 15.428 48.263 15.484 48.463 ;
 RECT 16.352 48.3635 16.408 48.5635 ;
 RECT 16.856 48.1115 16.912 48.3115 ;
 RECT 17.864 48.767 17.92 48.967 ;
 RECT 17.864 46.2015 17.92 46.4015 ;
 RECT 17.696 48.767 17.752 48.967 ;
 RECT 17.696 46.203 17.752 46.403 ;
 RECT 17.528 48.767 17.584 48.967 ;
 RECT 17.528 46.2015 17.584 46.4015 ;
 RECT 17.36 48.767 17.416 48.967 ;
 RECT 17.36 46.2015 17.416 46.4015 ;
 RECT 17.192 48.767 17.248 48.967 ;
 RECT 17.192 46.2015 17.248 46.4015 ;
 RECT 18.032 48.767 18.088 48.967 ;
 RECT 18.032 46.2015 18.088 46.4015 ;
 RECT 17.024 48.83 17.08 49.03 ;
 RECT 17.024 46.3155 17.08 46.5155 ;
 END
 END vss.gds3812
 PIN vss.gds3813
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.17 46.3635 25.23 46.5635 ;
 END
 END vss.gds3813
 PIN vss.gds3814
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.002 46.3635 25.062 46.5635 ;
 END
 END vss.gds3814
 PIN vss.gds3815
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.834 46.3635 24.894 46.5635 ;
 END
 END vss.gds3815
 PIN vss.gds3816
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.498 46.3635 24.558 46.5635 ;
 END
 END vss.gds3816
 PIN vss.gds3817
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.33 46.3635 24.39 46.5635 ;
 END
 END vss.gds3817
 PIN vss.gds3818
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.162 46.3635 24.222 46.5635 ;
 END
 END vss.gds3818
 PIN vss.gds3819
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.382 46.3635 20.442 46.5635 ;
 END
 END vss.gds3819
 PIN vss.gds3820
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.55 46.3635 20.61 46.5635 ;
 END
 END vss.gds3820
 PIN vss.gds3821
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.718 46.3635 20.778 46.5635 ;
 END
 END vss.gds3821
 PIN vss.gds3822
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.054 46.3635 21.114 46.5635 ;
 END
 END vss.gds3822
 PIN vss.gds3823
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.222 46.3635 21.282 46.5635 ;
 END
 END vss.gds3823
 PIN vss.gds3824
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.39 46.3635 21.45 46.5635 ;
 END
 END vss.gds3824
 PIN vss.gds3825
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.726 46.3635 21.786 46.5635 ;
 END
 END vss.gds3825
 PIN vss.gds3826
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.894 46.3635 21.954 46.5635 ;
 END
 END vss.gds3826
 PIN vss.gds3827
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.062 46.3635 22.122 46.5635 ;
 END
 END vss.gds3827
 PIN vss.gds3828
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 24.666 47.128 24.726 47.328 ;
 END
 END vss.gds3828
 PIN vss.gds3829
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 21.558 47.128 21.618 47.328 ;
 END
 END vss.gds3829
 PIN vss.gds3830
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 20.886 47.128 20.946 47.328 ;
 END
 END vss.gds3830
 PIN vss.gds3831
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.23 47.128 22.29 47.328 ;
 END
 END vss.gds3831
 PIN vss.gds3832
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.398 46.3635 22.458 46.5635 ;
 END
 END vss.gds3832
 PIN vss.gds3833
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.566 46.3635 22.626 46.5635 ;
 END
 END vss.gds3833
 PIN vss.gds3834
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.734 46.3635 22.794 46.5635 ;
 END
 END vss.gds3834
 PIN vss.gds3835
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.07 46.3635 23.13 46.5635 ;
 END
 END vss.gds3835
 PIN vss.gds3836
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.238 46.3635 23.298 46.5635 ;
 END
 END vss.gds3836
 PIN vss.gds3837
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.406 46.3635 23.466 46.5635 ;
 END
 END vss.gds3837
 PIN vss.gds3838
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 22.902 47.128 22.962 47.328 ;
 END
 END vss.gds3838
 PIN vss.gds3839
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 23.574 47.128 23.634 47.328 ;
 END
 END vss.gds3839
 PIN vss.gds3840
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 23.912 46.94 23.968 47.14 ;
 RECT 23.912 45.68 23.968 45.88 ;
 RECT 23.912 48.2 23.968 48.4 ;
 RECT 23.744 47.2135 23.8 47.4135 ;
 END
 END vss.gds3840
 PIN vss.gds3841
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.202 46.3635 29.262 46.5635 ;
 END
 END vss.gds3841
 PIN vss.gds3842
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.034 46.3635 29.094 46.5635 ;
 END
 END vss.gds3842
 PIN vss.gds3843
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.866 46.3635 28.926 46.5635 ;
 END
 END vss.gds3843
 PIN vss.gds3844
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.53 46.3635 28.59 46.5635 ;
 END
 END vss.gds3844
 PIN vss.gds3845
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.362 46.3635 28.422 46.5635 ;
 END
 END vss.gds3845
 PIN vss.gds3846
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.194 46.3635 28.254 46.5635 ;
 END
 END vss.gds3846
 PIN vss.gds3847
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.858 46.3635 27.918 46.5635 ;
 END
 END vss.gds3847
 PIN vss.gds3848
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.69 46.3635 27.75 46.5635 ;
 END
 END vss.gds3848
 PIN vss.gds3849
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.522 46.3635 27.582 46.5635 ;
 END
 END vss.gds3849
 PIN vss.gds3850
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.186 46.3635 27.246 46.5635 ;
 END
 END vss.gds3850
 PIN vss.gds3851
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.018 46.3635 27.078 46.5635 ;
 END
 END vss.gds3851
 PIN vss.gds3852
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.85 46.3635 26.91 46.5635 ;
 END
 END vss.gds3852
 PIN vss.gds3853
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.514 46.3635 26.574 46.5635 ;
 END
 END vss.gds3853
 PIN vss.gds3854
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.346 46.3635 26.406 46.5635 ;
 END
 END vss.gds3854
 PIN vss.gds3855
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.178 46.3635 26.238 46.5635 ;
 END
 END vss.gds3855
 PIN vss.gds3856
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.842 46.3635 25.902 46.5635 ;
 END
 END vss.gds3856
 PIN vss.gds3857
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.674 46.3635 25.734 46.5635 ;
 END
 END vss.gds3857
 PIN vss.gds3858
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.506 46.3635 25.566 46.5635 ;
 END
 END vss.gds3858
 PIN vss.gds3859
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.698 47.128 28.758 47.328 ;
 END
 END vss.gds3859
 PIN vss.gds3860
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 28.026 47.128 28.086 47.328 ;
 END
 END vss.gds3860
 PIN vss.gds3861
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 27.354 47.128 27.414 47.328 ;
 END
 END vss.gds3861
 PIN vss.gds3862
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.682 47.128 26.742 47.328 ;
 END
 END vss.gds3862
 PIN vss.gds3863
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 26.01 47.128 26.07 47.328 ;
 END
 END vss.gds3863
 PIN vss.gds3864
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 25.338 47.128 25.398 47.328 ;
 END
 END vss.gds3864
 PIN vss.gds3865
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.37 47.1405 29.43 47.3405 ;
 END
 END vss.gds3865
 PIN vss.gds3866
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.054 46.728 30.11 46.928 ;
 END
 END vss.gds3866
 PIN vss.gds3867
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.794 47.157 29.87 47.357 ;
 END
 END vss.gds3867
 PIN vss.gds3868
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 29.602 47.407 29.642 47.607 ;
 END
 END vss.gds3868
 PIN vss.gds3869
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 29.876 48.767 29.932 48.967 ;
 RECT 29.876 46.1645 29.932 46.3645 ;
 RECT 29.708 48.767 29.764 48.967 ;
 RECT 29.708 46.2015 29.764 46.4015 ;
 RECT 30.212 48.767 30.268 48.967 ;
 RECT 30.212 46.1645 30.268 46.3645 ;
 RECT 29.54 48.767 29.596 48.967 ;
 RECT 29.54 46.2015 29.596 46.4015 ;
 RECT 30.044 48.767 30.1 48.967 ;
 RECT 30.044 46.1645 30.1 46.3645 ;
 END
 END vss.gds3869
 PIN vss.gds3870
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 47.322 31.922 47.522 ;
 END
 END vss.gds3870
 PIN vss.gds3871
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 48.542 30.95 48.742 ;
 END
 END vss.gds3871
 PIN vss.gds3872
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 48.582 31.922 48.782 ;
 END
 END vss.gds3872
 PIN vss.gds3873
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.882 46.062 31.922 46.262 ;
 END
 END vss.gds3873
 PIN vss.gds3874
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 47.282 30.95 47.482 ;
 END
 END vss.gds3874
 PIN vss.gds3875
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.314 47.937 30.37 48.137 ;
 END
 END vss.gds3875
 PIN vss.gds3876
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.894 46.022 30.95 46.222 ;
 END
 END vss.gds3876
 PIN vss.gds3877
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.49 47.6795 34.546 47.8795 ;
 END
 END vss.gds3877
 PIN vss.gds3878
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 46.777 33.198 46.977 ;
 END
 END vss.gds3878
 PIN vss.gds3879
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.81 46.6495 33.866 46.8495 ;
 END
 END vss.gds3879
 PIN vss.gds3880
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 45.517 33.198 45.717 ;
 END
 END vss.gds3880
 PIN vss.gds3881
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.154 47.283 32.214 47.483 ;
 END
 END vss.gds3881
 PIN vss.gds3882
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.97 47.2205 34.046 47.4205 ;
 END
 END vss.gds3882
 PIN vss.gds3883
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.31 48.039 34.366 48.239 ;
 END
 END vss.gds3883
 PIN vss.gds3884
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.43 48.15 32.47 48.35 ;
 END
 END vss.gds3884
 PIN vss.gds3885
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.038 46.147 35.078 46.347 ;
 END
 END vss.gds3885
 PIN vss.gds3886
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 30.634 47.128 30.71 47.328 ;
 END
 END vss.gds3886
 PIN vss.gds3887
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 32.818 47.283 32.894 47.483 ;
 END
 END vss.gds3887
 PIN vss.gds3888
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.466 47.1965 33.542 47.3965 ;
 END
 END vss.gds3888
 PIN vss.gds3889
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 33.152 48.037 33.198 48.237 ;
 END
 END vss.gds3889
 PIN vss.gds3890
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 31.474 47.283 31.55 47.483 ;
 END
 END vss.gds3890
 PIN vss.gds3891
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 34.81 47.157 34.886 47.357 ;
 END
 END vss.gds3891
 PIN vss.gds3892
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 32.648 47.704 32.704 47.904 ;
 RECT 32.9 47.707 32.956 47.907 ;
 RECT 33.572 48.74 33.628 48.893 ;
 RECT 31.052 48.72 31.108 48.893 ;
 RECT 31.22 48.693 31.276 48.893 ;
 RECT 32.816 48.737 32.872 48.902 ;
 RECT 32.648 48.737 32.704 48.902 ;
 RECT 31.892 48.737 31.948 48.902 ;
 RECT 31.724 48.737 31.78 48.902 ;
 RECT 33.572 47.48 33.628 47.633 ;
 RECT 31.052 47.46 31.108 47.633 ;
 RECT 31.22 47.433 31.276 47.633 ;
 RECT 32.816 47.477 32.872 47.642 ;
 RECT 32.648 47.477 32.704 47.642 ;
 RECT 31.892 47.477 31.948 47.642 ;
 RECT 31.724 47.477 31.78 47.642 ;
 RECT 31.388 48.053 31.444 48.253 ;
 RECT 31.22 48.053 31.276 48.253 ;
 RECT 30.716 48.187 30.772 48.387 ;
 RECT 32.648 46.444 32.704 46.644 ;
 RECT 32.9 46.447 32.956 46.647 ;
 RECT 33.572 46.22 33.628 46.373 ;
 RECT 31.052 46.2 31.108 46.373 ;
 RECT 31.22 46.173 31.276 46.373 ;
 RECT 32.816 46.217 32.872 46.382 ;
 RECT 32.648 46.217 32.704 46.382 ;
 RECT 31.892 46.217 31.948 46.382 ;
 RECT 31.724 46.217 31.78 46.382 ;
 RECT 32.06 48.263 32.116 48.463 ;
 RECT 32.48 48.263 32.536 48.463 ;
 RECT 31.388 45.533 31.444 45.733 ;
 RECT 31.22 45.533 31.276 45.733 ;
 RECT 32.06 45.743 32.116 45.943 ;
 RECT 32.48 45.743 32.536 45.943 ;
 RECT 33.908 45.5915 33.964 45.7915 ;
 RECT 33.404 45.8435 33.46 46.0435 ;
 RECT 33.908 46.8515 33.964 47.0515 ;
 RECT 33.404 47.1035 33.46 47.3035 ;
 RECT 32.06 47.003 32.116 47.203 ;
 RECT 32.48 47.003 32.536 47.203 ;
 RECT 31.388 46.793 31.444 46.993 ;
 RECT 31.22 46.793 31.276 46.993 ;
 RECT 30.716 46.927 30.772 47.127 ;
 RECT 30.716 45.667 30.772 45.867 ;
 RECT 30.548 46.239 30.604 46.439 ;
 RECT 33.404 48.3635 33.46 48.5635 ;
 RECT 33.908 48.1115 33.964 48.3115 ;
 RECT 34.916 48.767 34.972 48.967 ;
 RECT 34.916 46.2015 34.972 46.4015 ;
 RECT 32.228 48.83 32.284 49.03 ;
 RECT 32.228 46.3665 32.284 46.5665 ;
 RECT 30.38 48.767 30.436 48.967 ;
 RECT 30.38 46.1045 30.436 46.3045 ;
 RECT 34.748 48.767 34.804 48.967 ;
 RECT 34.748 46.203 34.804 46.403 ;
 RECT 34.58 48.767 34.636 48.967 ;
 RECT 34.58 46.2015 34.636 46.4015 ;
 RECT 34.412 48.767 34.468 48.967 ;
 RECT 34.412 46.2015 34.468 46.4015 ;
 RECT 34.244 48.767 34.3 48.967 ;
 RECT 34.244 46.2015 34.3 46.4015 ;
 RECT 34.076 48.83 34.132 49.03 ;
 RECT 34.076 46.3155 34.132 46.5155 ;
 RECT 35.084 48.767 35.14 48.967 ;
 RECT 35.084 46.2015 35.14 46.4015 ;
 END
 END vss.gds3892
 PIN vss.gds3893
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.122 46.3635 40.182 46.5635 ;
 END
 END vss.gds3893
 PIN vss.gds3894
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.754 46.3635 35.814 46.5635 ;
 END
 END vss.gds3894
 PIN vss.gds3895
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.09 46.3635 36.15 46.5635 ;
 END
 END vss.gds3895
 PIN vss.gds3896
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.258 46.3635 36.318 46.5635 ;
 END
 END vss.gds3896
 PIN vss.gds3897
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.426 46.3635 36.486 46.5635 ;
 END
 END vss.gds3897
 PIN vss.gds3898
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.594 47.128 36.654 47.328 ;
 END
 END vss.gds3898
 PIN vss.gds3899
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.762 46.3635 36.822 46.5635 ;
 END
 END vss.gds3899
 PIN vss.gds3900
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 36.93 46.3635 36.99 46.5635 ;
 END
 END vss.gds3900
 PIN vss.gds3901
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.098 46.3635 37.158 46.5635 ;
 END
 END vss.gds3901
 PIN vss.gds3902
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.266 47.128 37.326 47.328 ;
 END
 END vss.gds3902
 PIN vss.gds3903
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.434 46.3635 37.494 46.5635 ;
 END
 END vss.gds3903
 PIN vss.gds3904
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.602 46.3635 37.662 46.5635 ;
 END
 END vss.gds3904
 PIN vss.gds3905
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.77 46.3635 37.83 46.5635 ;
 END
 END vss.gds3905
 PIN vss.gds3906
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 37.938 47.128 37.998 47.328 ;
 END
 END vss.gds3906
 PIN vss.gds3907
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.106 46.3635 38.166 46.5635 ;
 END
 END vss.gds3907
 PIN vss.gds3908
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.274 46.3635 38.334 46.5635 ;
 END
 END vss.gds3908
 PIN vss.gds3909
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.442 46.3635 38.502 46.5635 ;
 END
 END vss.gds3909
 PIN vss.gds3910
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.778 46.3635 38.838 46.5635 ;
 END
 END vss.gds3910
 PIN vss.gds3911
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.946 46.3635 39.006 46.5635 ;
 END
 END vss.gds3911
 PIN vss.gds3912
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.45 46.3635 39.51 46.5635 ;
 END
 END vss.gds3912
 PIN vss.gds3913
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.618 46.3635 39.678 46.5635 ;
 END
 END vss.gds3913
 PIN vss.gds3914
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.586 46.3635 35.646 46.5635 ;
 END
 END vss.gds3914
 PIN vss.gds3915
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.786 46.3635 39.846 46.5635 ;
 END
 END vss.gds3915
 PIN vss.gds3916
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.114 46.3635 39.174 46.5635 ;
 END
 END vss.gds3916
 PIN vss.gds3917
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.418 46.3635 35.478 46.5635 ;
 END
 END vss.gds3917
 PIN vss.gds3918
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 38.61 47.128 38.67 47.328 ;
 END
 END vss.gds3918
 PIN vss.gds3919
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.922 47.128 35.982 47.328 ;
 END
 END vss.gds3919
 PIN vss.gds3920
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.954 47.128 40.014 47.328 ;
 END
 END vss.gds3920
 PIN vss.gds3921
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 35.25 47.1405 35.31 47.3405 ;
 END
 END vss.gds3921
 PIN vss.gds3922
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 39.282 47.128 39.342 47.328 ;
 END
 END vss.gds3922
 PIN vss.gds3923
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.078 47.128 45.138 47.328 ;
 END
 END vss.gds3923
 PIN vss.gds3924
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.91 46.3635 44.97 46.5635 ;
 END
 END vss.gds3924
 PIN vss.gds3925
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.742 46.3635 44.802 46.5635 ;
 END
 END vss.gds3925
 PIN vss.gds3926
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.574 46.3635 44.634 46.5635 ;
 END
 END vss.gds3926
 PIN vss.gds3927
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.406 47.128 44.466 47.328 ;
 END
 END vss.gds3927
 PIN vss.gds3928
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.238 46.3635 44.298 46.5635 ;
 END
 END vss.gds3928
 PIN vss.gds3929
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 44.07 46.3635 44.13 46.5635 ;
 END
 END vss.gds3929
 PIN vss.gds3930
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.902 46.3635 43.962 46.5635 ;
 END
 END vss.gds3930
 PIN vss.gds3931
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.734 47.128 43.794 47.328 ;
 END
 END vss.gds3931
 PIN vss.gds3932
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.566 46.3635 43.626 46.5635 ;
 END
 END vss.gds3932
 PIN vss.gds3933
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.398 46.3635 43.458 46.5635 ;
 END
 END vss.gds3933
 PIN vss.gds3934
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.23 46.3635 43.29 46.5635 ;
 END
 END vss.gds3934
 PIN vss.gds3935
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 43.062 47.128 43.122 47.328 ;
 END
 END vss.gds3935
 PIN vss.gds3936
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.894 46.3635 42.954 46.5635 ;
 END
 END vss.gds3936
 PIN vss.gds3937
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.726 46.3635 42.786 46.5635 ;
 END
 END vss.gds3937
 PIN vss.gds3938
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.558 46.3635 42.618 46.5635 ;
 END
 END vss.gds3938
 PIN vss.gds3939
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.39 47.128 42.45 47.328 ;
 END
 END vss.gds3939
 PIN vss.gds3940
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.222 46.3635 42.282 46.5635 ;
 END
 END vss.gds3940
 PIN vss.gds3941
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 42.054 46.3635 42.114 46.5635 ;
 END
 END vss.gds3941
 PIN vss.gds3942
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.886 46.3635 41.946 46.5635 ;
 END
 END vss.gds3942
 PIN vss.gds3943
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.718 47.128 41.778 47.328 ;
 END
 END vss.gds3943
 PIN vss.gds3944
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.55 46.3635 41.61 46.5635 ;
 END
 END vss.gds3944
 PIN vss.gds3945
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.382 46.3635 41.442 46.5635 ;
 END
 END vss.gds3945
 PIN vss.gds3946
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 41.214 46.3635 41.274 46.5635 ;
 END
 END vss.gds3946
 PIN vss.gds3947
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.29 46.3635 40.35 46.5635 ;
 END
 END vss.gds3947
 PIN vss.gds3948
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.458 46.3635 40.518 46.5635 ;
 END
 END vss.gds3948
 PIN vss.gds3949
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 40.626 47.128 40.686 47.328 ;
 END
 END vss.gds3949
 PIN vss.gds3950
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 40.964 45.68 41.02 45.88 ;
 RECT 40.964 46.94 41.02 47.14 ;
 RECT 40.964 48.2 41.02 48.4 ;
 RECT 40.796 47.2135 40.852 47.4135 ;
 END
 END vss.gds3950
 PIN vss.gds3951
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 47.322 48.974 47.522 ;
 END
 END vss.gds3951
 PIN vss.gds3952
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 48.542 48.002 48.742 ;
 END
 END vss.gds3952
 PIN vss.gds3953
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 48.582 48.974 48.782 ;
 END
 END vss.gds3953
 PIN vss.gds3954
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.934 46.062 48.974 46.262 ;
 END
 END vss.gds3954
 PIN vss.gds3955
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 46.022 48.002 46.222 ;
 END
 END vss.gds3955
 PIN vss.gds3956
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.366 47.937 47.422 48.137 ;
 END
 END vss.gds3956
 PIN vss.gds3957
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.422 47.1405 46.482 47.3405 ;
 END
 END vss.gds3957
 PIN vss.gds3958
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.254 46.3635 46.314 46.5635 ;
 END
 END vss.gds3958
 PIN vss.gds3959
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.086 46.3635 46.146 46.5635 ;
 END
 END vss.gds3959
 PIN vss.gds3960
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.918 46.3635 45.978 46.5635 ;
 END
 END vss.gds3960
 PIN vss.gds3961
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.75 47.128 45.81 47.328 ;
 END
 END vss.gds3961
 PIN vss.gds3962
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.582 46.3635 45.642 46.5635 ;
 END
 END vss.gds3962
 PIN vss.gds3963
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.414 46.3635 45.474 46.5635 ;
 END
 END vss.gds3963
 PIN vss.gds3964
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 45.246 46.3635 45.306 46.5635 ;
 END
 END vss.gds3964
 PIN vss.gds3965
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.946 47.282 48.002 47.482 ;
 END
 END vss.gds3965
 PIN vss.gds3966
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 45.517 50.25 45.717 ;
 END
 END vss.gds3966
 PIN vss.gds3967
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 46.777 50.25 46.977 ;
 END
 END vss.gds3967
 PIN vss.gds3968
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.106 46.728 47.162 46.928 ;
 END
 END vss.gds3968
 PIN vss.gds3969
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.482 48.15 49.522 48.35 ;
 END
 END vss.gds3969
 PIN vss.gds3970
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.846 47.157 46.922 47.357 ;
 END
 END vss.gds3970
 PIN vss.gds3971
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 46.654 47.407 46.694 47.607 ;
 END
 END vss.gds3971
 PIN vss.gds3972
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 47.686 47.128 47.762 47.328 ;
 END
 END vss.gds3972
 PIN vss.gds3973
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.206 47.283 49.266 47.483 ;
 END
 END vss.gds3973
 PIN vss.gds3974
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 48.526 47.283 48.602 47.483 ;
 END
 END vss.gds3974
 PIN vss.gds3975
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 49.87 47.283 49.946 47.483 ;
 END
 END vss.gds3975
 PIN vss.gds3976
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.204 48.037 50.25 48.237 ;
 END
 END vss.gds3976
 PIN vss.gds3977
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 49.7 47.704 49.756 47.904 ;
 RECT 49.952 47.707 50.008 47.907 ;
 RECT 48.104 48.72 48.16 48.893 ;
 RECT 48.272 48.693 48.328 48.893 ;
 RECT 49.868 48.737 49.924 48.902 ;
 RECT 49.7 48.737 49.756 48.902 ;
 RECT 48.944 48.737 49 48.902 ;
 RECT 48.776 48.737 48.832 48.902 ;
 RECT 48.104 47.46 48.16 47.633 ;
 RECT 48.272 47.433 48.328 47.633 ;
 RECT 49.868 47.477 49.924 47.642 ;
 RECT 49.7 47.477 49.756 47.642 ;
 RECT 48.944 47.477 49 47.642 ;
 RECT 48.776 47.477 48.832 47.642 ;
 RECT 48.104 46.2 48.16 46.373 ;
 RECT 48.272 46.173 48.328 46.373 ;
 RECT 49.868 46.217 49.924 46.382 ;
 RECT 49.7 46.217 49.756 46.382 ;
 RECT 48.944 46.217 49 46.382 ;
 RECT 48.776 46.217 48.832 46.382 ;
 RECT 48.44 48.053 48.496 48.253 ;
 RECT 48.272 48.053 48.328 48.253 ;
 RECT 47.768 48.187 47.824 48.387 ;
 RECT 49.7 46.444 49.756 46.644 ;
 RECT 49.952 46.447 50.008 46.647 ;
 RECT 49.112 48.263 49.168 48.463 ;
 RECT 49.532 48.263 49.588 48.463 ;
 RECT 48.44 45.533 48.496 45.733 ;
 RECT 48.272 45.533 48.328 45.733 ;
 RECT 49.112 47.003 49.168 47.203 ;
 RECT 49.532 47.003 49.588 47.203 ;
 RECT 48.44 46.793 48.496 46.993 ;
 RECT 48.272 46.793 48.328 46.993 ;
 RECT 47.768 46.927 47.824 47.127 ;
 RECT 47.768 45.667 47.824 45.867 ;
 RECT 49.112 45.743 49.168 45.943 ;
 RECT 49.532 45.743 49.588 45.943 ;
 RECT 47.6 46.239 47.656 46.439 ;
 RECT 49.28 48.83 49.336 49.03 ;
 RECT 49.28 46.3665 49.336 46.5665 ;
 RECT 46.928 48.767 46.984 48.967 ;
 RECT 46.928 46.1645 46.984 46.3645 ;
 RECT 47.432 48.767 47.488 48.967 ;
 RECT 47.432 46.1045 47.488 46.3045 ;
 RECT 47.264 48.767 47.32 48.967 ;
 RECT 47.264 46.1645 47.32 46.3645 ;
 RECT 46.592 48.767 46.648 48.967 ;
 RECT 46.592 46.2015 46.648 46.4015 ;
 RECT 46.76 48.767 46.816 48.967 ;
 RECT 46.76 46.2015 46.816 46.4015 ;
 RECT 47.096 48.767 47.152 48.967 ;
 RECT 47.096 46.1645 47.152 46.3645 ;
 END
 END vss.gds3977
 PIN vss.gds3978
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.542 47.6795 51.598 47.8795 ;
 END
 END vss.gds3978
 PIN vss.gds3979
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.862 46.6495 50.918 46.8495 ;
 END
 END vss.gds3979
 PIN vss.gds3980
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.638 46.3635 52.698 46.5635 ;
 END
 END vss.gds3980
 PIN vss.gds3981
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.806 46.3635 52.866 46.5635 ;
 END
 END vss.gds3981
 PIN vss.gds3982
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.142 46.3635 53.202 46.5635 ;
 END
 END vss.gds3982
 PIN vss.gds3983
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.31 46.3635 53.37 46.5635 ;
 END
 END vss.gds3983
 PIN vss.gds3984
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.478 46.3635 53.538 46.5635 ;
 END
 END vss.gds3984
 PIN vss.gds3985
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.814 46.3635 53.874 46.5635 ;
 END
 END vss.gds3985
 PIN vss.gds3986
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.982 46.3635 54.042 46.5635 ;
 END
 END vss.gds3986
 PIN vss.gds3987
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.15 46.3635 54.21 46.5635 ;
 END
 END vss.gds3987
 PIN vss.gds3988
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.486 46.3635 54.546 46.5635 ;
 END
 END vss.gds3988
 PIN vss.gds3989
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.654 46.3635 54.714 46.5635 ;
 END
 END vss.gds3989
 PIN vss.gds3990
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.822 46.3635 54.882 46.5635 ;
 END
 END vss.gds3990
 PIN vss.gds3991
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.99 47.128 55.05 47.328 ;
 END
 END vss.gds3991
 PIN vss.gds3992
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.158 46.3635 55.218 46.5635 ;
 END
 END vss.gds3992
 PIN vss.gds3993
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 54.318 47.128 54.378 47.328 ;
 END
 END vss.gds3993
 PIN vss.gds3994
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 53.646 47.128 53.706 47.328 ;
 END
 END vss.gds3994
 PIN vss.gds3995
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.47 46.3635 52.53 46.5635 ;
 END
 END vss.gds3995
 PIN vss.gds3996
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.362 48.039 51.418 48.239 ;
 END
 END vss.gds3996
 PIN vss.gds3997
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.09 46.147 52.13 46.347 ;
 END
 END vss.gds3997
 PIN vss.gds3998
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.022 47.2205 51.098 47.4205 ;
 END
 END vss.gds3998
 PIN vss.gds3999
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.974 47.128 53.034 47.328 ;
 END
 END vss.gds3999
 PIN vss.gds4000
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 51.862 47.157 51.938 47.357 ;
 END
 END vss.gds4000
 PIN vss.gds4001
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 50.518 47.1965 50.594 47.3965 ;
 END
 END vss.gds4001
 PIN vss.gds4002
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 52.302 47.1405 52.362 47.3405 ;
 END
 END vss.gds4002
 PIN vss.gds4003
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 50.624 48.74 50.68 48.893 ;
 RECT 50.624 47.48 50.68 47.633 ;
 RECT 50.624 46.22 50.68 46.373 ;
 RECT 50.456 45.8435 50.512 46.0435 ;
 RECT 50.96 45.5915 51.016 45.7915 ;
 RECT 50.456 47.1035 50.512 47.3035 ;
 RECT 50.96 46.8515 51.016 47.0515 ;
 RECT 50.456 48.3635 50.512 48.5635 ;
 RECT 50.96 48.1115 51.016 48.3115 ;
 RECT 51.968 48.767 52.024 48.967 ;
 RECT 51.968 46.2015 52.024 46.4015 ;
 RECT 51.8 48.767 51.856 48.967 ;
 RECT 51.8 46.203 51.856 46.403 ;
 RECT 51.632 48.767 51.688 48.967 ;
 RECT 51.632 46.2015 51.688 46.4015 ;
 RECT 51.464 48.767 51.52 48.967 ;
 RECT 51.464 46.2015 51.52 46.4015 ;
 RECT 51.296 48.767 51.352 48.967 ;
 RECT 51.296 46.2015 51.352 46.4015 ;
 RECT 51.128 48.83 51.184 49.03 ;
 RECT 51.128 46.3155 51.184 46.5155 ;
 RECT 52.136 48.767 52.192 48.967 ;
 RECT 52.136 46.2015 52.192 46.4015 ;
 END
 END vss.gds4003
 PIN vss.gds4004
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.114 47.128 60.174 47.328 ;
 END
 END vss.gds4004
 PIN vss.gds4005
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.946 46.3635 60.006 46.5635 ;
 END
 END vss.gds4005
 PIN vss.gds4006
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.778 46.3635 59.838 46.5635 ;
 END
 END vss.gds4006
 PIN vss.gds4007
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.61 46.3635 59.67 46.5635 ;
 END
 END vss.gds4007
 PIN vss.gds4008
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.442 47.128 59.502 47.328 ;
 END
 END vss.gds4008
 PIN vss.gds4009
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.274 46.3635 59.334 46.5635 ;
 END
 END vss.gds4009
 PIN vss.gds4010
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 59.106 46.3635 59.166 46.5635 ;
 END
 END vss.gds4010
 PIN vss.gds4011
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.938 46.3635 58.998 46.5635 ;
 END
 END vss.gds4011
 PIN vss.gds4012
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.77 47.128 58.83 47.328 ;
 END
 END vss.gds4012
 PIN vss.gds4013
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.602 46.3635 58.662 46.5635 ;
 END
 END vss.gds4013
 PIN vss.gds4014
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.434 46.3635 58.494 46.5635 ;
 END
 END vss.gds4014
 PIN vss.gds4015
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 58.266 46.3635 58.326 46.5635 ;
 END
 END vss.gds4015
 PIN vss.gds4016
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.326 46.3635 55.386 46.5635 ;
 END
 END vss.gds4016
 PIN vss.gds4017
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.494 46.3635 55.554 46.5635 ;
 END
 END vss.gds4017
 PIN vss.gds4018
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.83 46.3635 55.89 46.5635 ;
 END
 END vss.gds4018
 PIN vss.gds4019
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.998 46.3635 56.058 46.5635 ;
 END
 END vss.gds4019
 PIN vss.gds4020
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.166 46.3635 56.226 46.5635 ;
 END
 END vss.gds4020
 PIN vss.gds4021
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.502 46.3635 56.562 46.5635 ;
 END
 END vss.gds4021
 PIN vss.gds4022
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.67 46.3635 56.73 46.5635 ;
 END
 END vss.gds4022
 PIN vss.gds4023
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.838 46.3635 56.898 46.5635 ;
 END
 END vss.gds4023
 PIN vss.gds4024
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.342 46.3635 57.402 46.5635 ;
 END
 END vss.gds4024
 PIN vss.gds4025
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.51 46.3635 57.57 46.5635 ;
 END
 END vss.gds4025
 PIN vss.gds4026
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 55.662 47.128 55.722 47.328 ;
 END
 END vss.gds4026
 PIN vss.gds4027
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 56.334 47.128 56.394 47.328 ;
 END
 END vss.gds4027
 PIN vss.gds4028
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.174 46.3635 57.234 46.5635 ;
 END
 END vss.gds4028
 PIN vss.gds4029
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.678 47.128 57.738 47.328 ;
 END
 END vss.gds4029
 PIN vss.gds4030
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 57.006 47.128 57.066 47.328 ;
 END
 END vss.gds4030
 PIN vss.gds4031
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 58.016 45.68 58.072 45.88 ;
 RECT 58.016 46.94 58.072 47.14 ;
 RECT 58.016 48.2 58.072 48.4 ;
 RECT 57.848 47.2135 57.904 47.4135 ;
 END
 END vss.gds4031
 PIN vss.gds4032
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 48.542 65.054 48.742 ;
 END
 END vss.gds4032
 PIN vss.gds4033
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.158 46.728 64.214 46.928 ;
 END
 END vss.gds4033
 PIN vss.gds4034
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.418 47.937 64.474 48.137 ;
 END
 END vss.gds4034
 PIN vss.gds4035
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.474 47.1405 63.534 47.3405 ;
 END
 END vss.gds4035
 PIN vss.gds4036
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.306 46.3635 63.366 46.5635 ;
 END
 END vss.gds4036
 PIN vss.gds4037
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.138 46.3635 63.198 46.5635 ;
 END
 END vss.gds4037
 PIN vss.gds4038
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.97 46.3635 63.03 46.5635 ;
 END
 END vss.gds4038
 PIN vss.gds4039
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.802 47.128 62.862 47.328 ;
 END
 END vss.gds4039
 PIN vss.gds4040
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.634 46.3635 62.694 46.5635 ;
 END
 END vss.gds4040
 PIN vss.gds4041
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.466 46.3635 62.526 46.5635 ;
 END
 END vss.gds4041
 PIN vss.gds4042
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.298 46.3635 62.358 46.5635 ;
 END
 END vss.gds4042
 PIN vss.gds4043
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 62.13 47.128 62.19 47.328 ;
 END
 END vss.gds4043
 PIN vss.gds4044
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.962 46.3635 62.022 46.5635 ;
 END
 END vss.gds4044
 PIN vss.gds4045
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.794 46.3635 61.854 46.5635 ;
 END
 END vss.gds4045
 PIN vss.gds4046
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.626 46.3635 61.686 46.5635 ;
 END
 END vss.gds4046
 PIN vss.gds4047
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.458 47.128 61.518 47.328 ;
 END
 END vss.gds4047
 PIN vss.gds4048
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.29 46.3635 61.35 46.5635 ;
 END
 END vss.gds4048
 PIN vss.gds4049
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 61.122 46.3635 61.182 46.5635 ;
 END
 END vss.gds4049
 PIN vss.gds4050
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.954 46.3635 61.014 46.5635 ;
 END
 END vss.gds4050
 PIN vss.gds4051
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.786 47.128 60.846 47.328 ;
 END
 END vss.gds4051
 PIN vss.gds4052
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.618 46.3635 60.678 46.5635 ;
 END
 END vss.gds4052
 PIN vss.gds4053
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.45 46.3635 60.51 46.5635 ;
 END
 END vss.gds4053
 PIN vss.gds4054
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 60.282 46.3635 60.342 46.5635 ;
 END
 END vss.gds4054
 PIN vss.gds4055
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.898 47.157 63.974 47.357 ;
 END
 END vss.gds4055
 PIN vss.gds4056
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 63.706 47.407 63.746 47.607 ;
 END
 END vss.gds4056
 PIN vss.gds4057
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 47.282 65.054 47.482 ;
 END
 END vss.gds4057
 PIN vss.gds4058
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.998 46.022 65.054 46.222 ;
 END
 END vss.gds4058
 PIN vss.gds4059
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 64.738 47.128 64.814 47.328 ;
 END
 END vss.gds4059
 PIN vss.gds4060
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 65.156 48.72 65.212 48.893 ;
 RECT 65.156 47.46 65.212 47.633 ;
 RECT 65.156 46.2 65.212 46.373 ;
 RECT 64.82 48.187 64.876 48.387 ;
 RECT 64.82 46.927 64.876 47.127 ;
 RECT 64.82 45.667 64.876 45.867 ;
 RECT 64.652 46.239 64.708 46.439 ;
 RECT 63.98 48.767 64.036 48.967 ;
 RECT 63.98 46.1645 64.036 46.3645 ;
 RECT 63.812 48.767 63.868 48.967 ;
 RECT 63.812 46.2015 63.868 46.4015 ;
 RECT 64.484 48.767 64.54 48.967 ;
 RECT 64.484 46.1045 64.54 46.3045 ;
 RECT 64.316 48.767 64.372 48.967 ;
 RECT 64.316 46.1645 64.372 46.3645 ;
 RECT 63.644 48.767 63.7 48.967 ;
 RECT 63.644 46.2015 63.7 46.4015 ;
 RECT 64.148 48.767 64.204 48.967 ;
 RECT 64.148 46.1645 64.204 46.3645 ;
 END
 END vss.gds4060
 PIN vss.gds4061
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 47.322 66.026 47.522 ;
 END
 END vss.gds4061
 PIN vss.gds4062
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 48.582 66.026 48.782 ;
 END
 END vss.gds4062
 PIN vss.gds4063
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.986 46.062 66.026 46.262 ;
 END
 END vss.gds4063
 PIN vss.gds4064
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 45.517 67.302 45.717 ;
 END
 END vss.gds4064
 PIN vss.gds4065
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.534 48.15 66.574 48.35 ;
 END
 END vss.gds4065
 PIN vss.gds4066
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.594 47.6795 68.65 47.8795 ;
 END
 END vss.gds4066
 PIN vss.gds4067
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 48.037 67.302 48.237 ;
 END
 END vss.gds4067
 PIN vss.gds4068
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.256 46.777 67.302 46.977 ;
 END
 END vss.gds4068
 PIN vss.gds4069
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.074 47.2205 68.15 47.4205 ;
 END
 END vss.gds4069
 PIN vss.gds4070
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.858 46.3635 69.918 46.5635 ;
 END
 END vss.gds4070
 PIN vss.gds4071
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.194 46.3635 70.254 46.5635 ;
 END
 END vss.gds4071
 PIN vss.gds4072
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.142 46.147 69.182 46.347 ;
 END
 END vss.gds4072
 PIN vss.gds4073
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.914 46.6495 67.97 46.8495 ;
 END
 END vss.gds4073
 PIN vss.gds4074
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.69 46.3635 69.75 46.5635 ;
 END
 END vss.gds4074
 PIN vss.gds4075
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.258 47.283 66.318 47.483 ;
 END
 END vss.gds4075
 PIN vss.gds4076
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.522 46.3635 69.582 46.5635 ;
 END
 END vss.gds4076
 PIN vss.gds4077
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.414 48.039 68.47 48.239 ;
 END
 END vss.gds4077
 PIN vss.gds4078
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.026 47.128 70.086 47.328 ;
 END
 END vss.gds4078
 PIN vss.gds4079
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 66.922 47.283 66.998 47.483 ;
 END
 END vss.gds4079
 PIN vss.gds4080
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 65.578 47.283 65.654 47.483 ;
 END
 END vss.gds4080
 PIN vss.gds4081
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 67.57 47.1965 67.646 47.3965 ;
 END
 END vss.gds4081
 PIN vss.gds4082
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 68.914 47.157 68.99 47.357 ;
 END
 END vss.gds4082
 PIN vss.gds4083
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 69.354 47.1405 69.414 47.3405 ;
 END
 END vss.gds4083
 PIN vss.gds4084
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m1 ;
 RECT 66.752 47.704 66.808 47.904 ;
 RECT 67.004 47.707 67.06 47.907 ;
 RECT 67.676 48.74 67.732 48.893 ;
 RECT 65.324 48.693 65.38 48.893 ;
 RECT 66.92 48.737 66.976 48.902 ;
 RECT 66.752 48.737 66.808 48.902 ;
 RECT 65.996 48.737 66.052 48.902 ;
 RECT 65.828 48.737 65.884 48.902 ;
 RECT 67.676 47.48 67.732 47.633 ;
 RECT 65.324 47.433 65.38 47.633 ;
 RECT 66.92 47.477 66.976 47.642 ;
 RECT 66.752 47.477 66.808 47.642 ;
 RECT 65.996 47.477 66.052 47.642 ;
 RECT 65.828 47.477 65.884 47.642 ;
 RECT 67.676 46.22 67.732 46.373 ;
 RECT 65.324 46.173 65.38 46.373 ;
 RECT 66.92 46.217 66.976 46.382 ;
 RECT 66.752 46.217 66.808 46.382 ;
 RECT 65.996 46.217 66.052 46.382 ;
 RECT 65.828 46.217 65.884 46.382 ;
 RECT 65.492 48.053 65.548 48.253 ;
 RECT 65.324 48.053 65.38 48.253 ;
 RECT 66.752 46.444 66.808 46.644 ;
 RECT 67.004 46.447 67.06 46.647 ;
 RECT 68.012 48.1115 68.068 48.3115 ;
 RECT 67.508 48.3635 67.564 48.5635 ;
 RECT 66.164 48.263 66.22 48.463 ;
 RECT 66.584 48.263 66.64 48.463 ;
 RECT 65.492 45.533 65.548 45.733 ;
 RECT 65.324 45.533 65.38 45.733 ;
 RECT 66.164 45.743 66.22 45.943 ;
 RECT 66.584 45.743 66.64 45.943 ;
 RECT 68.012 46.8515 68.068 47.0515 ;
 RECT 67.508 47.1035 67.564 47.3035 ;
 RECT 66.164 47.003 66.22 47.203 ;
 RECT 66.584 47.003 66.64 47.203 ;
 RECT 65.492 46.793 65.548 46.993 ;
 RECT 65.324 46.793 65.38 46.993 ;
 RECT 68.012 45.5915 68.068 45.7915 ;
 RECT 67.508 45.8435 67.564 46.0435 ;
 RECT 66.332 46.3665 66.388 46.5665 ;
 RECT 66.332 48.83 66.388 49.03 ;
 RECT 69.02 48.767 69.076 48.967 ;
 RECT 69.02 46.2015 69.076 46.4015 ;
 RECT 68.852 48.767 68.908 48.967 ;
 RECT 68.852 46.203 68.908 46.403 ;
 RECT 68.684 48.767 68.74 48.967 ;
 RECT 68.684 46.2015 68.74 46.4015 ;
 RECT 68.516 48.767 68.572 48.967 ;
 RECT 68.516 46.2015 68.572 46.4015 ;
 RECT 68.348 48.767 68.404 48.967 ;
 RECT 68.348 46.2015 68.404 46.4015 ;
 RECT 69.188 48.767 69.244 48.967 ;
 RECT 69.188 46.2015 69.244 46.4015 ;
 RECT 68.18 48.83 68.236 49.03 ;
 RECT 68.18 46.3155 68.236 46.5155 ;
 END
 END vss.gds4084
 PIN vss.gds4085
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.362 46.3635 70.422 46.5635 ;
 END
 END vss.gds4085
 PIN vss.gds4086
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.53 46.3635 70.59 46.5635 ;
 END
 END vss.gds4086
 PIN vss.gds4087
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.866 46.3635 70.926 46.5635 ;
 END
 END vss.gds4087
 PIN vss.gds4088
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.034 46.3635 71.094 46.5635 ;
 END
 END vss.gds4088
 PIN vss.gds4089
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.202 46.3635 71.262 46.5635 ;
 END
 END vss.gds4089
 PIN vss.gds4090
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.37 47.128 71.43 47.328 ;
 END
 END vss.gds4090
 PIN vss.gds4091
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.538 46.3635 71.598 46.5635 ;
 END
 END vss.gds4091
 PIN vss.gds4092
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.706 46.3635 71.766 46.5635 ;
 END
 END vss.gds4092
 PIN vss.gds4093
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 71.874 46.3635 71.934 46.5635 ;
 END
 END vss.gds4093
 PIN vss.gds4094
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.042 47.128 72.102 47.328 ;
 END
 END vss.gds4094
 PIN vss.gds4095
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.21 46.3635 72.27 46.5635 ;
 END
 END vss.gds4095
 PIN vss.gds4096
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.378 46.3635 72.438 46.5635 ;
 END
 END vss.gds4096
 PIN vss.gds4097
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.546 46.3635 72.606 46.5635 ;
 END
 END vss.gds4097
 PIN vss.gds4098
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.714 47.128 72.774 47.328 ;
 END
 END vss.gds4098
 PIN vss.gds4099
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 72.882 46.3635 72.942 46.5635 ;
 END
 END vss.gds4099
 PIN vss.gds4100
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.05 46.3635 73.11 46.5635 ;
 END
 END vss.gds4100
 PIN vss.gds4101
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.554 46.3635 73.614 46.5635 ;
 END
 END vss.gds4101
 PIN vss.gds4102
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.722 46.3635 73.782 46.5635 ;
 END
 END vss.gds4102
 PIN vss.gds4103
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.89 46.3635 73.95 46.5635 ;
 END
 END vss.gds4103
 PIN vss.gds4104
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.394 46.3635 74.454 46.5635 ;
 END
 END vss.gds4104
 PIN vss.gds4105
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.218 46.3635 73.278 46.5635 ;
 END
 END vss.gds4105
 PIN vss.gds4106
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.562 46.3635 74.622 46.5635 ;
 END
 END vss.gds4106
 PIN vss.gds4107
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.226 46.3635 74.286 46.5635 ;
 END
 END vss.gds4107
 PIN vss.gds4108
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 70.698 47.128 70.758 47.328 ;
 END
 END vss.gds4108
 PIN vss.gds4109
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 73.386 47.128 73.446 47.328 ;
 END
 END vss.gds4109
 PIN vss.gds4110
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.058 47.128 74.118 47.328 ;
 END
 END vss.gds4110
 PIN vss.gds4111
 DIRECTION INPUT ;
 USE GROUND ;
 PORT
 LAYER m3 ;
 RECT 74.73 47.128 74.79 47.328 ;
 END
 END vss.gds4111
 PIN vccdgt_1p0
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER m1 ;
 RECT 6.356 1.848 6.412 3.042 ;
 LAYER m1 ;
 RECT 6.356 3.108 6.412 4.302 ;
 LAYER m1 ;
 RECT 6.356 4.368 6.412 5.562 ;
 LAYER m1 ;
 RECT 6.356 5.628 6.412 6.822 ;
 LAYER m1 ;
 RECT 6.356 6.888 6.412 8.082 ;
 LAYER m1 ;
 RECT 6.356 8.148 6.412 9.342 ;
 LAYER m1 ;
 RECT 6.356 9.408 6.412 10.602 ;
 LAYER m1 ;
 RECT 6.356 10.668 6.412 11.862 ;
 LAYER m1 ;
 RECT 6.356 11.928 6.412 13.122 ;
 LAYER m1 ;
 RECT 6.356 13.188 6.412 14.382 ;
 LAYER m1 ;
 RECT 6.356 14.448 6.412 15.642 ;
 LAYER m1 ;
 RECT 6.356 15.708 6.412 16.902 ;
 LAYER m1 ;
 RECT 6.356 16.968 6.412 18.162 ;
 LAYER m1 ;
 RECT 6.356 18.228 6.412 19.422 ;
 LAYER m1 ;
 RECT 6.356 19.488 6.412 20.682 ;
 LAYER m1 ;
 RECT 7.532 28.464 7.588 28.532 ;
 LAYER m1 ;
 RECT 8.204 28.464 8.26 28.532 ;
 LAYER m1 ;
 RECT 8.876 28.464 8.932 28.532 ;
 LAYER m1 ;
 RECT 9.548 28.464 9.604 28.532 ;
 LAYER m1 ;
 RECT 10.22 28.464 10.276 28.532 ;
 LAYER m1 ;
 RECT 10.892 28.464 10.948 28.532 ;
 LAYER m1 ;
 RECT 11.564 28.464 11.62 28.532 ;
 LAYER m1 ;
 RECT 12.236 28.464 12.292 28.532 ;
 LAYER m1 ;
 RECT 18.788 28.464 18.844 28.532 ;
 LAYER m1 ;
 RECT 19.46 28.464 19.516 28.532 ;
 LAYER m1 ;
 RECT 17.192 28.602 17.248 28.672 ;
 LAYER m1 ;
 RECT 20.132 28.464 20.188 28.532 ;
 LAYER m1 ;
 RECT 20.804 28.464 20.86 28.532 ;
 LAYER m1 ;
 RECT 21.476 28.464 21.532 28.532 ;
 LAYER m1 ;
 RECT 22.148 28.464 22.204 28.532 ;
 LAYER m1 ;
 RECT 22.82 28.464 22.876 28.532 ;
 LAYER m1 ;
 RECT 23.492 28.464 23.548 28.532 ;
 LAYER m1 ;
 RECT 24.584 28.464 24.64 28.532 ;
 LAYER m1 ;
 RECT 25.256 28.464 25.312 28.532 ;
 LAYER m1 ;
 RECT 25.928 28.464 25.984 28.532 ;
 LAYER m1 ;
 RECT 26.6 28.464 26.656 28.532 ;
 LAYER m1 ;
 RECT 27.272 28.464 27.328 28.532 ;
 LAYER m1 ;
 RECT 27.944 28.464 28 28.532 ;
 LAYER m1 ;
 RECT 28.616 28.464 28.672 28.532 ;
 LAYER m1 ;
 RECT 29.288 28.464 29.344 28.532 ;
 LAYER m1 ;
 RECT 35.84 28.464 35.896 28.532 ;
 LAYER m1 ;
 RECT 36.512 28.464 36.568 28.532 ;
 LAYER m1 ;
 RECT 34.244 28.602 34.3 28.672 ;
 LAYER m1 ;
 RECT 37.184 28.464 37.24 28.532 ;
 LAYER m1 ;
 RECT 37.856 28.464 37.912 28.532 ;
 LAYER m1 ;
 RECT 38.528 28.464 38.584 28.532 ;
 LAYER m1 ;
 RECT 39.2 28.464 39.256 28.532 ;
 LAYER m1 ;
 RECT 39.872 28.464 39.928 28.532 ;
 LAYER m1 ;
 RECT 40.544 28.464 40.6 28.532 ;
 LAYER m1 ;
 RECT 41.636 28.464 41.692 28.532 ;
 LAYER m1 ;
 RECT 42.308 28.464 42.364 28.532 ;
 LAYER m1 ;
 RECT 42.98 28.464 43.036 28.532 ;
 LAYER m1 ;
 RECT 43.652 28.464 43.708 28.532 ;
 LAYER m1 ;
 RECT 44.324 28.464 44.38 28.532 ;
 LAYER m1 ;
 RECT 44.996 28.464 45.052 28.532 ;
 LAYER m1 ;
 RECT 45.668 28.464 45.724 28.532 ;
 LAYER m1 ;
 RECT 46.34 28.464 46.396 28.532 ;
 LAYER m1 ;
 RECT 52.892 28.464 52.948 28.532 ;
 LAYER m1 ;
 RECT 53.564 28.464 53.62 28.532 ;
 LAYER m1 ;
 RECT 51.296 28.602 51.352 28.672 ;
 LAYER m1 ;
 RECT 54.236 28.464 54.292 28.532 ;
 LAYER m1 ;
 RECT 54.908 28.464 54.964 28.532 ;
 LAYER m1 ;
 RECT 55.58 28.464 55.636 28.532 ;
 LAYER m1 ;
 RECT 56.252 28.464 56.308 28.532 ;
 LAYER m1 ;
 RECT 56.924 28.464 56.98 28.532 ;
 LAYER m1 ;
 RECT 57.596 28.464 57.652 28.532 ;
 LAYER m1 ;
 RECT 58.688 28.464 58.744 28.532 ;
 LAYER m1 ;
 RECT 59.36 28.464 59.416 28.532 ;
 LAYER m1 ;
 RECT 60.032 28.464 60.088 28.532 ;
 LAYER m1 ;
 RECT 60.704 28.464 60.76 28.532 ;
 LAYER m1 ;
 RECT 61.376 28.464 61.432 28.532 ;
 LAYER m1 ;
 RECT 62.048 28.464 62.104 28.532 ;
 LAYER m1 ;
 RECT 62.72 28.464 62.776 28.532 ;
 LAYER m1 ;
 RECT 63.392 28.464 63.448 28.532 ;
 LAYER m1 ;
 RECT 69.944 28.464 70 28.532 ;
 LAYER m1 ;
 RECT 70.616 28.464 70.672 28.532 ;
 LAYER m1 ;
 RECT 68.348 28.602 68.404 28.672 ;
 LAYER m1 ;
 RECT 71.288 28.464 71.344 28.532 ;
 LAYER m1 ;
 RECT 71.96 28.464 72.016 28.532 ;
 LAYER m1 ;
 RECT 72.632 28.464 72.688 28.532 ;
 LAYER m1 ;
 RECT 73.304 28.464 73.36 28.532 ;
 LAYER m1 ;
 RECT 73.976 28.464 74.032 28.532 ;
 LAYER m1 ;
 RECT 74.648 28.464 74.704 28.532 ;
 LAYER m1 ;
 RECT 6.356 28.812 6.412 30.006 ;
 LAYER m1 ;
 RECT 6.356 30.072 6.412 31.266 ;
 LAYER m1 ;
 RECT 6.356 31.332 6.412 32.526 ;
 LAYER m1 ;
 RECT 6.356 32.592 6.412 33.786 ;
 LAYER m1 ;
 RECT 6.356 33.852 6.412 35.046 ;
 LAYER m1 ;
 RECT 6.356 35.112 6.412 36.306 ;
 LAYER m1 ;
 RECT 6.356 36.372 6.412 37.566 ;
 LAYER m1 ;
 RECT 6.356 37.632 6.412 38.826 ;
 LAYER m1 ;
 RECT 6.356 38.892 6.412 40.086 ;
 LAYER m1 ;
 RECT 6.356 40.152 6.412 41.346 ;
 LAYER m1 ;
 RECT 6.356 41.412 6.412 42.606 ;
 LAYER m1 ;
 RECT 6.356 42.672 6.412 43.866 ;
 LAYER m1 ;
 RECT 6.356 43.932 6.412 45.126 ;
 LAYER m1 ;
 RECT 6.356 45.192 6.412 46.386 ;
 LAYER m1 ;
 RECT 6.356 46.452 6.412 47.646 ;
 LAYER m1 ;
 RECT 6.356 47.712 6.412 48.906 ;
 END
 END vccdgt_1p0
END c73p1rfshdxrom2048x32hb4img108_APACHECELL

END LIBRARY
