VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf104b064e1r1w0cbbehbaa4acw
  CLASS BLOCK ;
  FOREIGN arf104b064e1r1w0cbbehbaa4acw ;
  ORIGIN 0 0 ;
  SIZE 27 BY 24.96 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 13.8 14.316 15 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 11.88 11.528 13.08 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 13.8 15.516 15 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 13.8 10.028 15 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 13.8 10.116 15 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 13.8 10.372 15 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 13.8 10.628 15 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 13.8 10.716 15 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 13.8 14.528 15 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 13.8 14.616 15 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 13.8 14.872 15 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 13.8 15.128 15 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 11.88 12.816 13.08 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 11.88 13.072 13.08 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 11.88 13.328 13.08 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 11.88 13.416 13.08 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 11.88 13.628 13.08 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 11.88 14.228 13.08 ;
    END
  END wraddrp0[5]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 11.88 11.616 13.08 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 11.88 12.172 13.08 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 0.24 12.172 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 22.8 12.516 24 ;
    END
  END wrdatap0[100]
  PIN wrdatap0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 22.8 12.728 24 ;
    END
  END wrdatap0[101]
  PIN wrdatap0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 22.8 13.072 24 ;
    END
  END wrdatap0[102]
  PIN wrdatap0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 22.8 13.328 24 ;
    END
  END wrdatap0[103]
  PIN wrdatap0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 23.52 11.828 24.72 ;
    END
  END wrdatap0[104]
  PIN wrdatap0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 23.52 11.916 24.72 ;
    END
  END wrdatap0[105]
  PIN wrdatap0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 23.52 13.716 24.72 ;
    END
  END wrdatap0[106]
  PIN wrdatap0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 23.52 13.972 24.72 ;
    END
  END wrdatap0[107]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 1.68 13.716 2.88 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 1.68 13.972 2.88 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 2.4 12.516 3.6 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 2.4 12.728 3.6 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 2.4 13.072 3.6 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 2.4 13.328 3.6 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 3.12 11.828 4.32 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 3.12 11.916 4.32 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 3.12 13.716 4.32 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 3.12 13.972 4.32 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 0.24 12.428 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 3.84 12.516 5.04 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 3.84 12.728 5.04 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 3.84 13.072 5.04 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 3.84 13.328 5.04 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 4.56 11.828 5.76 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 4.56 11.916 5.76 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 4.56 13.716 5.76 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 4.56 13.972 5.76 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 5.28 12.516 6.48 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 5.28 12.728 6.48 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 0.24 13.716 1.44 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 5.28 13.072 6.48 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 5.28 13.328 6.48 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 6 11.828 7.2 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 6 11.916 7.2 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 6 13.716 7.2 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 6 13.972 7.2 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 6.72 12.516 7.92 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 6.72 12.728 7.92 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 6.72 13.072 7.92 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 6.72 13.328 7.92 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 0.24 13.972 1.44 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 7.44 11.828 8.64 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 7.44 11.916 8.64 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 7.44 13.716 8.64 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 7.44 13.972 8.64 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 8.16 12.516 9.36 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 8.16 12.728 9.36 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 8.16 13.072 9.36 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 8.16 13.328 9.36 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 8.88 11.828 10.08 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 8.88 11.916 10.08 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 0.96 12.516 2.16 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 8.88 13.716 10.08 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 8.88 13.972 10.08 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 9.6 12.516 10.8 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 9.6 12.728 10.8 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 9.6 13.072 10.8 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 9.6 13.328 10.8 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 10.32 11.828 11.52 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 10.32 11.916 11.52 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 10.32 13.716 11.52 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 10.32 13.972 11.52 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 0.96 12.728 2.16 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 15.6 12.172 16.8 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 15.6 12.428 16.8 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 15.6 13.716 16.8 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 15.6 13.972 16.8 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 16.32 12.816 17.52 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 16.32 11.828 17.52 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 16.32 13.328 17.52 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 16.32 13.416 17.52 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 17.04 12.172 18.24 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 17.04 12.428 18.24 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 0.96 13.072 2.16 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 17.04 13.972 18.24 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 17.04 13.072 18.24 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 17.76 11.828 18.96 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 17.76 11.916 18.96 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 17.76 13.628 18.96 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 17.76 13.716 18.96 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 18.48 12.516 19.68 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 18.48 12.728 19.68 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 18.48 13.072 19.68 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 18.48 13.328 19.68 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 0.96 13.328 2.16 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 19.2 11.828 20.4 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 19.2 11.916 20.4 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 19.2 13.716 20.4 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 19.2 13.972 20.4 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 19.92 12.516 21.12 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 19.92 12.728 21.12 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 19.92 13.072 21.12 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 19.92 13.328 21.12 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 20.64 11.828 21.84 ;
    END
  END wrdatap0[88]
  PIN wrdatap0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 20.64 11.916 21.84 ;
    END
  END wrdatap0[89]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 1.68 11.828 2.88 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 20.64 13.716 21.84 ;
    END
  END wrdatap0[90]
  PIN wrdatap0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 20.64 13.972 21.84 ;
    END
  END wrdatap0[91]
  PIN wrdatap0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 21.36 12.516 22.56 ;
    END
  END wrdatap0[92]
  PIN wrdatap0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 21.36 12.728 22.56 ;
    END
  END wrdatap0[93]
  PIN wrdatap0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 21.36 13.072 22.56 ;
    END
  END wrdatap0[94]
  PIN wrdatap0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 21.36 13.328 22.56 ;
    END
  END wrdatap0[95]
  PIN wrdatap0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 22.08 11.828 23.28 ;
    END
  END wrdatap0[96]
  PIN wrdatap0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 22.08 11.916 23.28 ;
    END
  END wrdatap0[97]
  PIN wrdatap0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 22.08 13.716 23.28 ;
    END
  END wrdatap0[98]
  PIN wrdatap0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 22.08 13.972 23.28 ;
    END
  END wrdatap0[99]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 1.68 11.916 2.88 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 11.88 12.516 13.08 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 11.88 12.728 13.08 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 11.88 12.428 13.08 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 0.24 10.028 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 22.8 10.028 24 ;
    END
  END rddatap0[100]
  PIN rddatap0[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 22.8 10.116 24 ;
    END
  END rddatap0[101]
  PIN rddatap0[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 22.8 14.528 24 ;
    END
  END rddatap0[102]
  PIN rddatap0[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 22.8 14.616 24 ;
    END
  END rddatap0[103]
  PIN rddatap0[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 23.52 11.016 24.72 ;
    END
  END rddatap0[104]
  PIN rddatap0[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 23.52 11.272 24.72 ;
    END
  END rddatap0[105]
  PIN rddatap0[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 23.52 15.216 24.72 ;
    END
  END rddatap0[106]
  PIN rddatap0[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 23.52 15.428 24.72 ;
    END
  END rddatap0[107]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 1.68 15.216 2.88 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 1.68 15.428 2.88 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 2.4 10.028 3.6 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 2.4 10.116 3.6 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 2.4 14.528 3.6 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 2.4 14.616 3.6 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 3.12 11.016 4.32 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 3.12 11.272 4.32 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 3.12 15.216 4.32 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 3.12 15.428 4.32 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 0.24 10.116 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 3.84 10.028 5.04 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 3.84 10.116 5.04 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 3.84 14.528 5.04 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 3.84 14.616 5.04 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 4.56 11.016 5.76 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 4.56 11.272 5.76 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 4.56 15.216 5.76 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 4.56 15.428 5.76 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 5.28 10.028 6.48 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 5.28 10.116 6.48 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 0.24 15.216 1.44 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 5.28 14.528 6.48 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 5.28 14.616 6.48 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 6 11.016 7.2 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 6 11.272 7.2 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 6 15.216 7.2 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 6 15.428 7.2 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 6.72 10.028 7.92 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 6.72 10.116 7.92 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 6.72 14.528 7.92 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 6.72 14.616 7.92 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 0.24 15.428 1.44 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 7.44 11.016 8.64 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 7.44 11.272 8.64 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 7.44 15.216 8.64 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 7.44 15.428 8.64 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 8.16 10.028 9.36 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 8.16 10.116 9.36 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 8.16 14.528 9.36 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 8.16 14.616 9.36 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 8.88 11.016 10.08 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 8.88 11.272 10.08 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 0.96 10.372 2.16 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 8.88 15.216 10.08 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 8.88 15.428 10.08 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 9.6 10.028 10.8 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 9.6 10.116 10.8 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 9.6 14.528 10.8 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 9.6 14.616 10.8 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 10.32 11.016 11.52 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 10.32 11.272 11.52 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 10.32 15.216 11.52 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 10.32 15.428 11.52 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 0.96 10.628 2.16 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 15.6 10.928 16.8 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 15.6 11.016 16.8 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 15.6 14.228 16.8 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 15.6 15.216 16.8 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 16.32 10.372 17.52 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 16.32 10.628 17.52 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 16.32 14.872 17.52 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 16.32 15.128 17.52 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 17.04 11.272 18.24 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 17.04 10.028 18.24 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 0.96 14.528 2.16 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 17.04 14.316 18.24 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 17.04 14.528 18.24 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 17.76 10.716 18.96 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 17.76 10.928 18.96 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 17.76 15.216 18.96 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 17.76 15.428 18.96 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 18.48 10.028 19.68 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 18.48 10.116 19.68 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 18.48 14.528 19.68 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 18.48 14.616 19.68 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 0.96 14.616 2.16 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 19.2 11.016 20.4 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 19.2 11.272 20.4 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 19.2 15.216 20.4 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 19.2 15.428 20.4 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 19.92 10.028 21.12 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 19.92 10.116 21.12 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 19.92 14.528 21.12 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 19.92 14.616 21.12 ;
    END
  END rddatap0[87]
  PIN rddatap0[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 20.64 11.016 21.84 ;
    END
  END rddatap0[88]
  PIN rddatap0[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 20.64 11.272 21.84 ;
    END
  END rddatap0[89]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 1.68 11.016 2.88 ;
    END
  END rddatap0[8]
  PIN rddatap0[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 20.64 15.216 21.84 ;
    END
  END rddatap0[90]
  PIN rddatap0[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 20.64 15.428 21.84 ;
    END
  END rddatap0[91]
  PIN rddatap0[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 21.36 10.028 22.56 ;
    END
  END rddatap0[92]
  PIN rddatap0[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 21.36 10.116 22.56 ;
    END
  END rddatap0[93]
  PIN rddatap0[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 21.36 14.528 22.56 ;
    END
  END rddatap0[94]
  PIN rddatap0[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 21.36 14.616 22.56 ;
    END
  END rddatap0[95]
  PIN rddatap0[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 22.08 11.016 23.28 ;
    END
  END rddatap0[96]
  PIN rddatap0[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 22.08 11.272 23.28 ;
    END
  END rddatap0[97]
  PIN rddatap0[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 22.08 15.216 23.28 ;
    END
  END rddatap0[98]
  PIN rddatap0[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 22.08 15.428 23.28 ;
    END
  END rddatap0[99]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 1.68 11.272 2.88 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 24.9 ;
        RECT 2.662 0.06 2.738 24.9 ;
        RECT 4.462 0.06 4.538 24.9 ;
        RECT 6.262 0.06 6.338 24.9 ;
        RECT 8.062 0.06 8.138 24.9 ;
        RECT 9.862 0.06 9.938 24.9 ;
        RECT 11.662 0.06 11.738 24.9 ;
        RECT 13.462 0.06 13.538 24.9 ;
        RECT 15.262 0.06 15.338 24.9 ;
        RECT 17.062 0.06 17.138 24.9 ;
        RECT 18.862 0.06 18.938 24.9 ;
        RECT 20.662 0.06 20.738 24.9 ;
        RECT 22.462 0.06 22.538 24.9 ;
        RECT 24.262 0.06 24.338 24.9 ;
        RECT 26.062 0.06 26.138 24.9 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 24.9 ;
        RECT 3.562 0.06 3.638 24.9 ;
        RECT 5.362 0.06 5.438 24.9 ;
        RECT 7.162 0.06 7.238 24.9 ;
        RECT 8.962 0.06 9.038 24.9 ;
        RECT 10.762 0.06 10.838 24.9 ;
        RECT 12.562 0.06 12.638 24.9 ;
        RECT 14.362 0.06 14.438 24.9 ;
        RECT 16.162 0.06 16.238 24.9 ;
        RECT 17.962 0.06 18.038 24.9 ;
        RECT 19.762 0.06 19.838 24.9 ;
        RECT 21.562 0.06 21.638 24.9 ;
        RECT 23.362 0.06 23.438 24.9 ;
        RECT 25.162 0.06 25.238 24.9 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 27.016 24.974 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 27.02 24.98 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 27.0705 24.998 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 27.035 25.03 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 27.07 24.998 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 27.059 25.05 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 27.09 25.022 ;
    LAYER m7 SPACING 0 ;
      RECT 26.138 25.02 27.04 25.08 ;
      RECT 26.138 -0.06 27.092 25.02 ;
      RECT 26.138 -0.12 27.04 -0.06 ;
      RECT 25.238 -0.12 26.062 25.08 ;
      RECT 24.338 -0.12 25.162 25.08 ;
      RECT 23.438 -0.12 24.262 25.08 ;
      RECT 22.538 -0.12 23.362 25.08 ;
      RECT 21.638 -0.12 22.462 25.08 ;
      RECT 20.738 -0.12 21.562 25.08 ;
      RECT 19.838 -0.12 20.662 25.08 ;
      RECT 18.938 -0.12 19.762 25.08 ;
      RECT 18.038 -0.12 18.862 25.08 ;
      RECT 17.138 -0.12 17.962 25.08 ;
      RECT 16.238 -0.12 17.062 25.08 ;
      RECT 15.338 24.72 16.162 25.08 ;
      RECT 15.338 23.52 15.384 24.72 ;
      RECT 15.428 23.52 16.162 24.72 ;
      RECT 15.338 23.28 16.162 23.52 ;
      RECT 15.338 22.08 15.384 23.28 ;
      RECT 15.428 22.08 16.162 23.28 ;
      RECT 15.338 21.84 16.162 22.08 ;
      RECT 15.338 20.64 15.384 21.84 ;
      RECT 15.428 20.64 16.162 21.84 ;
      RECT 15.338 20.4 16.162 20.64 ;
      RECT 15.338 19.2 15.384 20.4 ;
      RECT 15.428 19.2 16.162 20.4 ;
      RECT 15.338 18.96 16.162 19.2 ;
      RECT 15.338 17.76 15.384 18.96 ;
      RECT 15.428 17.76 16.162 18.96 ;
      RECT 15.338 15 16.162 17.76 ;
      RECT 15.338 13.8 15.472 15 ;
      RECT 15.516 13.8 16.162 15 ;
      RECT 15.338 11.52 16.162 13.8 ;
      RECT 15.338 10.32 15.384 11.52 ;
      RECT 15.428 10.32 16.162 11.52 ;
      RECT 15.338 10.08 16.162 10.32 ;
      RECT 15.338 8.88 15.384 10.08 ;
      RECT 15.428 8.88 16.162 10.08 ;
      RECT 15.338 8.64 16.162 8.88 ;
      RECT 15.338 7.44 15.384 8.64 ;
      RECT 15.428 7.44 16.162 8.64 ;
      RECT 15.338 7.2 16.162 7.44 ;
      RECT 15.338 6 15.384 7.2 ;
      RECT 15.428 6 16.162 7.2 ;
      RECT 15.338 5.76 16.162 6 ;
      RECT 15.338 4.56 15.384 5.76 ;
      RECT 15.428 4.56 16.162 5.76 ;
      RECT 15.338 4.32 16.162 4.56 ;
      RECT 15.338 3.12 15.384 4.32 ;
      RECT 15.428 3.12 16.162 4.32 ;
      RECT 15.338 2.88 16.162 3.12 ;
      RECT 15.338 1.68 15.384 2.88 ;
      RECT 15.428 1.68 16.162 2.88 ;
      RECT 15.338 1.44 16.162 1.68 ;
      RECT 15.338 0.24 15.384 1.44 ;
      RECT 15.428 0.24 16.162 1.44 ;
      RECT 15.338 -0.12 16.162 0.24 ;
      RECT 14.438 24.72 15.262 25.08 ;
      RECT 14.438 24 15.172 24.72 ;
      RECT 15.216 23.52 15.262 24.72 ;
      RECT 14.616 23.52 15.172 24 ;
      RECT 14.616 23.28 15.262 23.52 ;
      RECT 14.438 22.8 14.484 24 ;
      RECT 14.528 22.8 14.572 24 ;
      RECT 14.616 22.8 15.172 23.28 ;
      RECT 14.438 22.56 15.172 22.8 ;
      RECT 15.216 22.08 15.262 23.28 ;
      RECT 14.616 22.08 15.172 22.56 ;
      RECT 14.616 21.84 15.262 22.08 ;
      RECT 14.438 21.36 14.484 22.56 ;
      RECT 14.528 21.36 14.572 22.56 ;
      RECT 14.616 21.36 15.172 21.84 ;
      RECT 14.438 21.12 15.172 21.36 ;
      RECT 15.216 20.64 15.262 21.84 ;
      RECT 14.616 20.64 15.172 21.12 ;
      RECT 14.616 20.4 15.262 20.64 ;
      RECT 14.438 19.92 14.484 21.12 ;
      RECT 14.528 19.92 14.572 21.12 ;
      RECT 14.616 19.92 15.172 20.4 ;
      RECT 14.438 19.68 15.172 19.92 ;
      RECT 15.216 19.2 15.262 20.4 ;
      RECT 14.616 19.2 15.172 19.68 ;
      RECT 14.616 18.96 15.262 19.2 ;
      RECT 14.438 18.48 14.484 19.68 ;
      RECT 14.528 18.48 14.572 19.68 ;
      RECT 14.616 18.48 15.172 18.96 ;
      RECT 14.438 18.24 15.172 18.48 ;
      RECT 15.216 17.76 15.262 18.96 ;
      RECT 14.528 17.76 15.172 18.24 ;
      RECT 14.528 17.52 15.262 17.76 ;
      RECT 14.438 17.04 14.484 18.24 ;
      RECT 14.528 17.04 14.828 17.52 ;
      RECT 15.128 16.8 15.262 17.52 ;
      RECT 14.872 16.32 15.084 17.52 ;
      RECT 14.438 16.32 14.828 17.04 ;
      RECT 15.128 16.32 15.172 16.8 ;
      RECT 15.216 15.6 15.262 16.8 ;
      RECT 14.438 15.6 15.172 16.32 ;
      RECT 14.438 15 15.262 15.6 ;
      RECT 14.438 13.8 14.484 15 ;
      RECT 14.528 13.8 14.572 15 ;
      RECT 14.616 13.8 14.828 15 ;
      RECT 14.872 13.8 15.084 15 ;
      RECT 15.128 13.8 15.262 15 ;
      RECT 14.438 11.52 15.262 13.8 ;
      RECT 14.438 10.8 15.172 11.52 ;
      RECT 15.216 10.32 15.262 11.52 ;
      RECT 14.616 10.32 15.172 10.8 ;
      RECT 14.616 10.08 15.262 10.32 ;
      RECT 14.438 9.6 14.484 10.8 ;
      RECT 14.528 9.6 14.572 10.8 ;
      RECT 14.616 9.6 15.172 10.08 ;
      RECT 14.438 9.36 15.172 9.6 ;
      RECT 15.216 8.88 15.262 10.08 ;
      RECT 14.616 8.88 15.172 9.36 ;
      RECT 14.616 8.64 15.262 8.88 ;
      RECT 14.438 8.16 14.484 9.36 ;
      RECT 14.528 8.16 14.572 9.36 ;
      RECT 14.616 8.16 15.172 8.64 ;
      RECT 14.438 7.92 15.172 8.16 ;
      RECT 15.216 7.44 15.262 8.64 ;
      RECT 14.616 7.44 15.172 7.92 ;
      RECT 14.616 7.2 15.262 7.44 ;
      RECT 14.438 6.72 14.484 7.92 ;
      RECT 14.528 6.72 14.572 7.92 ;
      RECT 14.616 6.72 15.172 7.2 ;
      RECT 14.438 6.48 15.172 6.72 ;
      RECT 15.216 6 15.262 7.2 ;
      RECT 14.616 6 15.172 6.48 ;
      RECT 14.616 5.76 15.262 6 ;
      RECT 14.438 5.28 14.484 6.48 ;
      RECT 14.528 5.28 14.572 6.48 ;
      RECT 14.616 5.28 15.172 5.76 ;
      RECT 14.438 5.04 15.172 5.28 ;
      RECT 15.216 4.56 15.262 5.76 ;
      RECT 14.616 4.56 15.172 5.04 ;
      RECT 14.616 4.32 15.262 4.56 ;
      RECT 14.438 3.84 14.484 5.04 ;
      RECT 14.528 3.84 14.572 5.04 ;
      RECT 14.616 3.84 15.172 4.32 ;
      RECT 14.438 3.6 15.172 3.84 ;
      RECT 15.216 3.12 15.262 4.32 ;
      RECT 14.616 3.12 15.172 3.6 ;
      RECT 14.616 2.88 15.262 3.12 ;
      RECT 14.438 2.4 14.484 3.6 ;
      RECT 14.528 2.4 14.572 3.6 ;
      RECT 14.616 2.4 15.172 2.88 ;
      RECT 14.438 2.16 15.172 2.4 ;
      RECT 15.216 1.68 15.262 2.88 ;
      RECT 14.616 1.68 15.172 2.16 ;
      RECT 14.616 1.44 15.262 1.68 ;
      RECT 14.438 0.96 14.484 2.16 ;
      RECT 14.528 0.96 14.572 2.16 ;
      RECT 14.616 0.96 15.172 1.44 ;
      RECT 15.216 0.24 15.262 1.44 ;
      RECT 14.438 0.24 15.172 0.96 ;
      RECT 14.438 -0.12 15.262 0.24 ;
      RECT 13.538 24.72 14.362 25.08 ;
      RECT 13.538 23.52 13.672 24.72 ;
      RECT 13.716 23.52 13.928 24.72 ;
      RECT 13.972 23.52 14.362 24.72 ;
      RECT 13.538 23.28 14.362 23.52 ;
      RECT 13.538 22.08 13.672 23.28 ;
      RECT 13.716 22.08 13.928 23.28 ;
      RECT 13.972 22.08 14.362 23.28 ;
      RECT 13.538 21.84 14.362 22.08 ;
      RECT 13.538 20.64 13.672 21.84 ;
      RECT 13.716 20.64 13.928 21.84 ;
      RECT 13.972 20.64 14.362 21.84 ;
      RECT 13.538 20.4 14.362 20.64 ;
      RECT 13.538 19.2 13.672 20.4 ;
      RECT 13.716 19.2 13.928 20.4 ;
      RECT 13.972 19.2 14.362 20.4 ;
      RECT 13.538 18.96 14.362 19.2 ;
      RECT 13.716 18.24 14.362 18.96 ;
      RECT 13.538 17.76 13.584 18.96 ;
      RECT 13.628 17.76 13.672 18.96 ;
      RECT 13.716 17.76 13.928 18.24 ;
      RECT 13.972 17.04 14.272 18.24 ;
      RECT 14.316 17.04 14.362 18.24 ;
      RECT 13.538 17.04 13.928 17.76 ;
      RECT 13.538 16.8 14.362 17.04 ;
      RECT 13.538 15.6 13.672 16.8 ;
      RECT 13.716 15.6 13.928 16.8 ;
      RECT 13.972 15.6 14.184 16.8 ;
      RECT 14.228 15.6 14.362 16.8 ;
      RECT 13.538 15 14.362 15.6 ;
      RECT 13.538 13.8 14.272 15 ;
      RECT 14.316 13.8 14.362 15 ;
      RECT 13.538 13.08 14.362 13.8 ;
      RECT 13.538 11.88 13.584 13.08 ;
      RECT 13.628 11.88 14.184 13.08 ;
      RECT 14.228 11.88 14.362 13.08 ;
      RECT 13.538 11.52 14.362 11.88 ;
      RECT 13.538 10.32 13.672 11.52 ;
      RECT 13.716 10.32 13.928 11.52 ;
      RECT 13.972 10.32 14.362 11.52 ;
      RECT 13.538 10.08 14.362 10.32 ;
      RECT 13.538 8.88 13.672 10.08 ;
      RECT 13.716 8.88 13.928 10.08 ;
      RECT 13.972 8.88 14.362 10.08 ;
      RECT 13.538 8.64 14.362 8.88 ;
      RECT 13.538 7.44 13.672 8.64 ;
      RECT 13.716 7.44 13.928 8.64 ;
      RECT 13.972 7.44 14.362 8.64 ;
      RECT 13.538 7.2 14.362 7.44 ;
      RECT 13.538 6 13.672 7.2 ;
      RECT 13.716 6 13.928 7.2 ;
      RECT 13.972 6 14.362 7.2 ;
      RECT 13.538 5.76 14.362 6 ;
      RECT 13.538 4.56 13.672 5.76 ;
      RECT 13.716 4.56 13.928 5.76 ;
      RECT 13.972 4.56 14.362 5.76 ;
      RECT 13.538 4.32 14.362 4.56 ;
      RECT 13.538 3.12 13.672 4.32 ;
      RECT 13.716 3.12 13.928 4.32 ;
      RECT 13.972 3.12 14.362 4.32 ;
      RECT 13.538 2.88 14.362 3.12 ;
      RECT 13.538 1.68 13.672 2.88 ;
      RECT 13.716 1.68 13.928 2.88 ;
      RECT 13.972 1.68 14.362 2.88 ;
      RECT 13.538 1.44 14.362 1.68 ;
      RECT 13.538 0.24 13.672 1.44 ;
      RECT 13.716 0.24 13.928 1.44 ;
      RECT 13.972 0.24 14.362 1.44 ;
      RECT 13.538 -0.12 14.362 0.24 ;
      RECT 12.638 24 13.462 25.08 ;
      RECT 12.638 22.8 12.684 24 ;
      RECT 12.728 22.8 13.028 24 ;
      RECT 13.072 22.8 13.284 24 ;
      RECT 13.328 22.8 13.462 24 ;
      RECT 12.638 22.56 13.462 22.8 ;
      RECT 12.638 21.36 12.684 22.56 ;
      RECT 12.728 21.36 13.028 22.56 ;
      RECT 13.072 21.36 13.284 22.56 ;
      RECT 13.328 21.36 13.462 22.56 ;
      RECT 12.638 21.12 13.462 21.36 ;
      RECT 12.638 19.92 12.684 21.12 ;
      RECT 12.728 19.92 13.028 21.12 ;
      RECT 13.072 19.92 13.284 21.12 ;
      RECT 13.328 19.92 13.462 21.12 ;
      RECT 12.638 19.68 13.462 19.92 ;
      RECT 12.638 18.48 12.684 19.68 ;
      RECT 12.728 18.48 13.028 19.68 ;
      RECT 13.072 18.48 13.284 19.68 ;
      RECT 13.328 18.48 13.462 19.68 ;
      RECT 12.638 18.24 13.462 18.48 ;
      RECT 12.638 17.52 13.028 18.24 ;
      RECT 13.072 17.52 13.462 18.24 ;
      RECT 12.816 17.04 13.028 17.52 ;
      RECT 13.072 17.04 13.284 17.52 ;
      RECT 12.638 16.32 12.772 17.52 ;
      RECT 13.328 16.32 13.372 17.52 ;
      RECT 13.416 16.32 13.462 17.52 ;
      RECT 12.816 16.32 13.284 17.04 ;
      RECT 12.638 13.08 13.462 16.32 ;
      RECT 12.638 11.88 12.684 13.08 ;
      RECT 12.728 11.88 12.772 13.08 ;
      RECT 12.816 11.88 13.028 13.08 ;
      RECT 13.072 11.88 13.284 13.08 ;
      RECT 13.328 11.88 13.372 13.08 ;
      RECT 13.416 11.88 13.462 13.08 ;
      RECT 12.638 10.8 13.462 11.88 ;
      RECT 12.638 9.6 12.684 10.8 ;
      RECT 12.728 9.6 13.028 10.8 ;
      RECT 13.072 9.6 13.284 10.8 ;
      RECT 13.328 9.6 13.462 10.8 ;
      RECT 12.638 9.36 13.462 9.6 ;
      RECT 12.638 8.16 12.684 9.36 ;
      RECT 12.728 8.16 13.028 9.36 ;
      RECT 13.072 8.16 13.284 9.36 ;
      RECT 13.328 8.16 13.462 9.36 ;
      RECT 12.638 7.92 13.462 8.16 ;
      RECT 12.638 6.72 12.684 7.92 ;
      RECT 12.728 6.72 13.028 7.92 ;
      RECT 13.072 6.72 13.284 7.92 ;
      RECT 13.328 6.72 13.462 7.92 ;
      RECT 12.638 6.48 13.462 6.72 ;
      RECT 12.638 5.28 12.684 6.48 ;
      RECT 12.728 5.28 13.028 6.48 ;
      RECT 13.072 5.28 13.284 6.48 ;
      RECT 13.328 5.28 13.462 6.48 ;
      RECT 12.638 5.04 13.462 5.28 ;
      RECT 12.638 3.84 12.684 5.04 ;
      RECT 12.728 3.84 13.028 5.04 ;
      RECT 13.072 3.84 13.284 5.04 ;
      RECT 13.328 3.84 13.462 5.04 ;
      RECT 12.638 3.6 13.462 3.84 ;
      RECT 12.638 2.4 12.684 3.6 ;
      RECT 12.728 2.4 13.028 3.6 ;
      RECT 13.072 2.4 13.284 3.6 ;
      RECT 13.328 2.4 13.462 3.6 ;
      RECT 12.638 2.16 13.462 2.4 ;
      RECT 12.638 0.96 12.684 2.16 ;
      RECT 12.728 0.96 13.028 2.16 ;
      RECT 13.072 0.96 13.284 2.16 ;
      RECT 13.328 0.96 13.462 2.16 ;
      RECT 12.638 -0.12 13.462 0.96 ;
      RECT 11.738 24.72 12.562 25.08 ;
      RECT 11.916 24 12.562 24.72 ;
      RECT 11.738 23.52 11.784 24.72 ;
      RECT 11.828 23.52 11.872 24.72 ;
      RECT 11.916 23.52 12.472 24 ;
      RECT 11.738 23.28 12.472 23.52 ;
      RECT 12.516 22.8 12.562 24 ;
      RECT 11.916 22.8 12.472 23.28 ;
      RECT 11.916 22.56 12.562 22.8 ;
      RECT 11.738 22.08 11.784 23.28 ;
      RECT 11.828 22.08 11.872 23.28 ;
      RECT 11.916 22.08 12.472 22.56 ;
      RECT 11.738 21.84 12.472 22.08 ;
      RECT 12.516 21.36 12.562 22.56 ;
      RECT 11.916 21.36 12.472 21.84 ;
      RECT 11.916 21.12 12.562 21.36 ;
      RECT 11.738 20.64 11.784 21.84 ;
      RECT 11.828 20.64 11.872 21.84 ;
      RECT 11.916 20.64 12.472 21.12 ;
      RECT 11.738 20.4 12.472 20.64 ;
      RECT 12.516 19.92 12.562 21.12 ;
      RECT 11.916 19.92 12.472 20.4 ;
      RECT 11.916 19.68 12.562 19.92 ;
      RECT 11.738 19.2 11.784 20.4 ;
      RECT 11.828 19.2 11.872 20.4 ;
      RECT 11.916 19.2 12.472 19.68 ;
      RECT 11.738 18.96 12.472 19.2 ;
      RECT 12.516 18.48 12.562 19.68 ;
      RECT 11.916 18.48 12.472 18.96 ;
      RECT 11.916 18.24 12.562 18.48 ;
      RECT 11.738 17.76 11.784 18.96 ;
      RECT 11.828 17.76 11.872 18.96 ;
      RECT 11.916 17.76 12.128 18.24 ;
      RECT 11.738 17.52 12.128 17.76 ;
      RECT 12.172 17.04 12.384 18.24 ;
      RECT 12.428 17.04 12.562 18.24 ;
      RECT 11.828 17.04 12.128 17.52 ;
      RECT 11.828 16.8 12.562 17.04 ;
      RECT 11.738 16.32 11.784 17.52 ;
      RECT 11.828 16.32 12.128 16.8 ;
      RECT 12.172 15.6 12.384 16.8 ;
      RECT 12.428 15.6 12.562 16.8 ;
      RECT 11.738 15.6 12.128 16.32 ;
      RECT 11.738 13.08 12.562 15.6 ;
      RECT 11.738 11.88 12.128 13.08 ;
      RECT 12.172 11.88 12.384 13.08 ;
      RECT 12.428 11.88 12.472 13.08 ;
      RECT 12.516 11.88 12.562 13.08 ;
      RECT 11.738 11.52 12.562 11.88 ;
      RECT 11.916 10.8 12.562 11.52 ;
      RECT 11.738 10.32 11.784 11.52 ;
      RECT 11.828 10.32 11.872 11.52 ;
      RECT 11.916 10.32 12.472 10.8 ;
      RECT 11.738 10.08 12.472 10.32 ;
      RECT 12.516 9.6 12.562 10.8 ;
      RECT 11.916 9.6 12.472 10.08 ;
      RECT 11.916 9.36 12.562 9.6 ;
      RECT 11.738 8.88 11.784 10.08 ;
      RECT 11.828 8.88 11.872 10.08 ;
      RECT 11.916 8.88 12.472 9.36 ;
      RECT 11.738 8.64 12.472 8.88 ;
      RECT 12.516 8.16 12.562 9.36 ;
      RECT 11.916 8.16 12.472 8.64 ;
      RECT 11.916 7.92 12.562 8.16 ;
      RECT 11.738 7.44 11.784 8.64 ;
      RECT 11.828 7.44 11.872 8.64 ;
      RECT 11.916 7.44 12.472 7.92 ;
      RECT 11.738 7.2 12.472 7.44 ;
      RECT 12.516 6.72 12.562 7.92 ;
      RECT 11.916 6.72 12.472 7.2 ;
      RECT 11.916 6.48 12.562 6.72 ;
      RECT 11.738 6 11.784 7.2 ;
      RECT 11.828 6 11.872 7.2 ;
      RECT 11.916 6 12.472 6.48 ;
      RECT 11.738 5.76 12.472 6 ;
      RECT 12.516 5.28 12.562 6.48 ;
      RECT 11.916 5.28 12.472 5.76 ;
      RECT 11.916 5.04 12.562 5.28 ;
      RECT 11.738 4.56 11.784 5.76 ;
      RECT 11.828 4.56 11.872 5.76 ;
      RECT 11.916 4.56 12.472 5.04 ;
      RECT 11.738 4.32 12.472 4.56 ;
      RECT 12.516 3.84 12.562 5.04 ;
      RECT 11.916 3.84 12.472 4.32 ;
      RECT 11.916 3.6 12.562 3.84 ;
      RECT 11.738 3.12 11.784 4.32 ;
      RECT 11.828 3.12 11.872 4.32 ;
      RECT 11.916 3.12 12.472 3.6 ;
      RECT 11.738 2.88 12.472 3.12 ;
      RECT 12.516 2.4 12.562 3.6 ;
      RECT 11.916 2.4 12.472 2.88 ;
      RECT 11.916 2.16 12.562 2.4 ;
      RECT 11.738 1.68 11.784 2.88 ;
      RECT 11.828 1.68 11.872 2.88 ;
      RECT 11.916 1.68 12.472 2.16 ;
      RECT 11.738 1.44 12.472 1.68 ;
      RECT 12.516 0.96 12.562 2.16 ;
      RECT 12.428 0.96 12.472 1.44 ;
      RECT 11.738 0.24 12.128 1.44 ;
      RECT 12.172 0.24 12.384 1.44 ;
      RECT 12.428 0.24 12.562 0.96 ;
      RECT 11.738 -0.12 12.562 0.24 ;
      RECT 10.838 24.72 11.662 25.08 ;
      RECT 10.838 23.52 10.972 24.72 ;
      RECT 11.016 23.52 11.228 24.72 ;
      RECT 11.272 23.52 11.662 24.72 ;
      RECT 10.838 23.28 11.662 23.52 ;
      RECT 10.838 22.08 10.972 23.28 ;
      RECT 11.016 22.08 11.228 23.28 ;
      RECT 11.272 22.08 11.662 23.28 ;
      RECT 10.838 21.84 11.662 22.08 ;
      RECT 10.838 20.64 10.972 21.84 ;
      RECT 11.016 20.64 11.228 21.84 ;
      RECT 11.272 20.64 11.662 21.84 ;
      RECT 10.838 20.4 11.662 20.64 ;
      RECT 10.838 19.2 10.972 20.4 ;
      RECT 11.016 19.2 11.228 20.4 ;
      RECT 11.272 19.2 11.662 20.4 ;
      RECT 10.838 18.96 11.662 19.2 ;
      RECT 10.928 18.24 11.662 18.96 ;
      RECT 10.838 17.76 10.884 18.96 ;
      RECT 10.928 17.76 11.228 18.24 ;
      RECT 11.272 17.04 11.662 18.24 ;
      RECT 10.838 17.04 11.228 17.76 ;
      RECT 10.838 16.8 11.662 17.04 ;
      RECT 10.838 15.6 10.884 16.8 ;
      RECT 10.928 15.6 10.972 16.8 ;
      RECT 11.016 15.6 11.662 16.8 ;
      RECT 10.838 13.08 11.662 15.6 ;
      RECT 10.838 11.88 11.484 13.08 ;
      RECT 11.528 11.88 11.572 13.08 ;
      RECT 11.616 11.88 11.662 13.08 ;
      RECT 10.838 11.52 11.662 11.88 ;
      RECT 10.838 10.32 10.972 11.52 ;
      RECT 11.016 10.32 11.228 11.52 ;
      RECT 11.272 10.32 11.662 11.52 ;
      RECT 10.838 10.08 11.662 10.32 ;
      RECT 10.838 8.88 10.972 10.08 ;
      RECT 11.016 8.88 11.228 10.08 ;
      RECT 11.272 8.88 11.662 10.08 ;
      RECT 10.838 8.64 11.662 8.88 ;
      RECT 10.838 7.44 10.972 8.64 ;
      RECT 11.016 7.44 11.228 8.64 ;
      RECT 11.272 7.44 11.662 8.64 ;
      RECT 10.838 7.2 11.662 7.44 ;
      RECT 10.838 6 10.972 7.2 ;
      RECT 11.016 6 11.228 7.2 ;
      RECT 11.272 6 11.662 7.2 ;
      RECT 10.838 5.76 11.662 6 ;
      RECT 10.838 4.56 10.972 5.76 ;
      RECT 11.016 4.56 11.228 5.76 ;
      RECT 11.272 4.56 11.662 5.76 ;
      RECT 10.838 4.32 11.662 4.56 ;
      RECT 10.838 3.12 10.972 4.32 ;
      RECT 11.016 3.12 11.228 4.32 ;
      RECT 11.272 3.12 11.662 4.32 ;
      RECT 10.838 2.88 11.662 3.12 ;
      RECT 10.838 1.68 10.972 2.88 ;
      RECT 11.016 1.68 11.228 2.88 ;
      RECT 11.272 1.68 11.662 2.88 ;
      RECT 10.838 -0.12 11.662 1.68 ;
      RECT 9.938 24 10.762 25.08 ;
      RECT 9.938 22.8 9.984 24 ;
      RECT 10.028 22.8 10.072 24 ;
      RECT 10.116 22.8 10.762 24 ;
      RECT 9.938 22.56 10.762 22.8 ;
      RECT 9.938 21.36 9.984 22.56 ;
      RECT 10.028 21.36 10.072 22.56 ;
      RECT 10.116 21.36 10.762 22.56 ;
      RECT 9.938 21.12 10.762 21.36 ;
      RECT 9.938 19.92 9.984 21.12 ;
      RECT 10.028 19.92 10.072 21.12 ;
      RECT 10.116 19.92 10.762 21.12 ;
      RECT 9.938 19.68 10.762 19.92 ;
      RECT 10.116 18.96 10.762 19.68 ;
      RECT 9.938 18.48 9.984 19.68 ;
      RECT 10.028 18.48 10.072 19.68 ;
      RECT 10.116 18.48 10.672 18.96 ;
      RECT 9.938 18.24 10.672 18.48 ;
      RECT 10.716 17.76 10.762 18.96 ;
      RECT 10.028 17.76 10.672 18.24 ;
      RECT 10.028 17.52 10.762 17.76 ;
      RECT 9.938 17.04 9.984 18.24 ;
      RECT 10.028 17.04 10.328 17.52 ;
      RECT 10.372 16.32 10.584 17.52 ;
      RECT 10.628 16.32 10.762 17.52 ;
      RECT 9.938 16.32 10.328 17.04 ;
      RECT 9.938 15 10.762 16.32 ;
      RECT 9.938 13.8 9.984 15 ;
      RECT 10.028 13.8 10.072 15 ;
      RECT 10.116 13.8 10.328 15 ;
      RECT 10.372 13.8 10.584 15 ;
      RECT 10.628 13.8 10.672 15 ;
      RECT 10.716 13.8 10.762 15 ;
      RECT 9.938 10.8 10.762 13.8 ;
      RECT 9.938 9.6 9.984 10.8 ;
      RECT 10.028 9.6 10.072 10.8 ;
      RECT 10.116 9.6 10.762 10.8 ;
      RECT 9.938 9.36 10.762 9.6 ;
      RECT 9.938 8.16 9.984 9.36 ;
      RECT 10.028 8.16 10.072 9.36 ;
      RECT 10.116 8.16 10.762 9.36 ;
      RECT 9.938 7.92 10.762 8.16 ;
      RECT 9.938 6.72 9.984 7.92 ;
      RECT 10.028 6.72 10.072 7.92 ;
      RECT 10.116 6.72 10.762 7.92 ;
      RECT 9.938 6.48 10.762 6.72 ;
      RECT 9.938 5.28 9.984 6.48 ;
      RECT 10.028 5.28 10.072 6.48 ;
      RECT 10.116 5.28 10.762 6.48 ;
      RECT 9.938 5.04 10.762 5.28 ;
      RECT 9.938 3.84 9.984 5.04 ;
      RECT 10.028 3.84 10.072 5.04 ;
      RECT 10.116 3.84 10.762 5.04 ;
      RECT 9.938 3.6 10.762 3.84 ;
      RECT 9.938 2.4 9.984 3.6 ;
      RECT 10.028 2.4 10.072 3.6 ;
      RECT 10.116 2.4 10.762 3.6 ;
      RECT 9.938 2.16 10.762 2.4 ;
      RECT 9.938 1.44 10.328 2.16 ;
      RECT 10.372 0.96 10.584 2.16 ;
      RECT 10.628 0.96 10.762 2.16 ;
      RECT 10.116 0.96 10.328 1.44 ;
      RECT 9.938 0.24 9.984 1.44 ;
      RECT 10.028 0.24 10.072 1.44 ;
      RECT 10.116 0.24 10.762 0.96 ;
      RECT 9.938 -0.12 10.762 0.24 ;
      RECT 9.038 -0.12 9.862 25.08 ;
      RECT 8.138 -0.12 8.962 25.08 ;
      RECT 7.238 -0.12 8.062 25.08 ;
      RECT 6.338 -0.12 7.162 25.08 ;
      RECT 5.438 -0.12 6.262 25.08 ;
      RECT 4.538 -0.12 5.362 25.08 ;
      RECT 3.638 -0.12 4.462 25.08 ;
      RECT 2.738 -0.12 3.562 25.08 ;
      RECT 1.838 -0.12 2.662 25.08 ;
      RECT 0.938 -0.12 1.762 25.08 ;
      RECT -0.04 25.02 0.862 25.08 ;
      RECT -0.092 -0.06 0.862 25.02 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 26.258 0 26.92 24.96 ;
      RECT 25.358 0 25.942 24.96 ;
      RECT 24.458 0 25.042 24.96 ;
      RECT 23.558 0 24.142 24.96 ;
      RECT 22.658 0 23.242 24.96 ;
      RECT 21.758 0 22.342 24.96 ;
      RECT 20.858 0 21.442 24.96 ;
      RECT 19.958 0 20.542 24.96 ;
      RECT 19.058 0 19.642 24.96 ;
      RECT 18.158 0 18.742 24.96 ;
      RECT 17.258 0 17.842 24.96 ;
      RECT 16.358 0 16.942 24.96 ;
      RECT 15.458 24.84 16.042 24.96 ;
      RECT 15.548 17.64 16.042 24.84 ;
      RECT 15.458 15.12 16.042 17.64 ;
      RECT 15.636 13.68 16.042 15.12 ;
      RECT 15.458 11.64 16.042 13.68 ;
      RECT 15.548 0.12 16.042 11.64 ;
      RECT 15.458 0 16.042 0.12 ;
      RECT 14.558 24.84 15.142 24.96 ;
      RECT 14.558 24.12 15.052 24.84 ;
      RECT 14.736 18.36 15.052 24.12 ;
      RECT 14.648 17.64 15.052 18.36 ;
      RECT 14.648 16.92 14.708 17.64 ;
      RECT 14.558 16.2 14.708 16.92 ;
      RECT 14.558 15.48 15.052 16.2 ;
      RECT 14.558 15.12 15.142 15.48 ;
      RECT 13.658 24.84 14.242 24.96 ;
      RECT 14.092 19.08 14.242 24.84 ;
      RECT 13.836 18.36 14.242 19.08 ;
      RECT 14.092 16.92 14.152 18.36 ;
      RECT 12.758 24.12 13.342 24.96 ;
      RECT 12.848 18.36 12.908 24.12 ;
      RECT 12.758 17.64 12.908 18.36 ;
      RECT 11.858 24.84 12.442 24.96 ;
      RECT 12.036 24.12 12.442 24.84 ;
      RECT 12.036 18.36 12.352 24.12 ;
      RECT 10.958 24.84 11.542 24.96 ;
      RECT 11.392 19.08 11.542 24.84 ;
      RECT 11.048 18.36 11.542 19.08 ;
      RECT 11.048 17.64 11.108 18.36 ;
      RECT 11.392 16.92 11.542 18.36 ;
      RECT 10.958 16.92 11.108 17.64 ;
      RECT 11.136 15.48 11.542 16.92 ;
      RECT 10.958 13.2 11.542 15.48 ;
      RECT 10.958 11.76 11.364 13.2 ;
      RECT 10.958 11.64 11.542 11.76 ;
      RECT 11.392 1.56 11.542 11.64 ;
      RECT 10.958 0 11.542 1.56 ;
      RECT 10.058 24.12 10.642 24.96 ;
      RECT 10.236 19.08 10.642 24.12 ;
      RECT 10.236 18.36 10.552 19.08 ;
      RECT 10.148 17.64 10.552 18.36 ;
      RECT 10.148 16.92 10.208 17.64 ;
      RECT 10.058 16.2 10.208 16.92 ;
      RECT 10.058 15.12 10.642 16.2 ;
      RECT 9.158 0 9.742 24.96 ;
      RECT 8.258 0 8.842 24.96 ;
      RECT 7.358 0 7.942 24.96 ;
      RECT 6.458 0 7.042 24.96 ;
      RECT 5.558 0 6.142 24.96 ;
      RECT 4.658 0 5.242 24.96 ;
      RECT 3.758 0 4.342 24.96 ;
      RECT 2.858 0 3.442 24.96 ;
      RECT 1.958 0 2.542 24.96 ;
      RECT 1.058 0 1.642 24.96 ;
      RECT 0.08 0 0.742 24.96 ;
      RECT 13.192 17.64 13.342 18.36 ;
      RECT 13.658 16.92 13.808 17.64 ;
      RECT 11.948 16.2 12.008 17.64 ;
      RECT 11.858 15.48 12.008 16.2 ;
      RECT 11.858 13.2 12.442 15.48 ;
      RECT 11.858 11.76 12.008 13.2 ;
      RECT 11.858 11.64 12.442 11.76 ;
      RECT 12.036 10.92 12.442 11.64 ;
      RECT 12.036 1.56 12.352 10.92 ;
      RECT 12.936 16.2 13.164 16.92 ;
      RECT 12.758 13.2 13.342 16.2 ;
      RECT 13.658 15.12 14.242 15.48 ;
      RECT 13.658 13.68 14.152 15.12 ;
      RECT 13.658 13.2 14.242 13.68 ;
      RECT 13.748 11.76 14.064 13.2 ;
      RECT 13.658 11.64 14.242 11.76 ;
      RECT 14.092 0.12 14.242 11.64 ;
      RECT 13.658 0 14.242 0.12 ;
      RECT 14.558 11.64 15.142 13.68 ;
      RECT 14.558 10.92 15.052 11.64 ;
      RECT 14.736 0.84 15.052 10.92 ;
      RECT 14.558 0.12 15.052 0.84 ;
      RECT 14.558 0 15.142 0.12 ;
      RECT 10.058 10.92 10.642 13.68 ;
      RECT 10.236 2.28 10.642 10.92 ;
      RECT 12.758 10.92 13.342 11.76 ;
      RECT 12.848 0.84 12.908 10.92 ;
      RECT 12.758 0 13.342 0.84 ;
      RECT 10.058 1.56 10.208 2.28 ;
      RECT 11.858 0.12 12.008 1.56 ;
      RECT 11.858 0 12.442 0.12 ;
      RECT 10.236 0.12 10.642 0.84 ;
      RECT 10.058 0 10.642 0.12 ;
    LAYER m0 ;
      RECT 0 0.002 27 24.958 ;
    LAYER m1 ;
      RECT 0 0 27 24.96 ;
    LAYER m2 ;
      RECT 0 0.015 27 24.945 ;
    LAYER m3 ;
      RECT 0.015 0 26.985 24.96 ;
    LAYER m4 ;
      RECT 0 0.02 27 24.94 ;
    LAYER m5 ;
      RECT 0.012 0 26.988 24.96 ;
    LAYER m6 ;
      RECT 0 0.012 27 24.948 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf104b064e1r1w0cbbehbaa4acw

END LIBRARY
