//-----------------------------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2020 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to the source code
// ("Material") are owned by Intel Corporation or its suppliers or licensors. Title to the Material
// remains with Intel Corporation or its suppliers and licensors. The Material contains trade
// secrets and proprietary and confidential information of Intel or its suppliers and licensors.
// The Material is protected by worldwide copyright and trade secret laws and treaty provisions.
// No part of the Material may be used, copied, reproduced, modified, published, uploaded, posted,
// transmitted, distributed, or disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual property right is
// granted to or conferred upon you by disclosure or delivery of the Materials, either expressly, by
// implication, inducement, estoppel or otherwise. Any license under such intellectual property rights
// must be express and approved by Intel in writing.
//
//-----------------------------------------------------------------------------------------------------
// AW_clkgate
//
// This module is responsible for implementing a 2-input clock "AND" gate w/ a latch on the enable.
//
//-----------------------------------------------------------------------------------------------------

module hqm_AW_clkgate (

     input  logic       clk                 // Input clock
    ,input  logic       enable              // Clock enable
    ,input  logic       cfg_clkungate       // CFG override to force ungating the clock
    ,input  logic       fscan_clkungate     // DFX override to force ungating the clock

    ,output logic       gated_clk           // Gated output clock
);

//-----------------------------------------------------------------------------------------------------

// collage-pragma translate_on

logic local_enable;

assign local_enable = enable | cfg_clkungate;

hqm_AW_ctech_clk_gate_te i_clkgate (

     .clk       (clk)
    ,.en        (local_enable)
    ,.te        (fscan_clkungate)
    ,.clkout    (gated_clk)
);

// collage-pragma translate_on

endmodule // AW_clkgate

