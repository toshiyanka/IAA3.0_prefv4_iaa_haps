class PowerGating;



	typedef enum {
		RST_ASD,
		RST_DSD,		
		SW_PG_REQ,
		DEASSERT_SW_PG_REQ,
		SW_PG_REQ_DSD,		
		//RESTORE commands
		SIP_RESTORE,
		DEASSERT_SIP_RESTORE,
		SIP_RESTORE_DSD,
		SIP_RESTORE_NEXT_WAKE,
		//RESTORE commands
		SIP_PG_ACK,
		SIP_UG_ACK,

		PMC_SIP_WAKE,
		DEASSERT_PMC_SIP_WAKE,		
		PMC_SIP_WAKE_DSD,

		FAB_PG_REQ,
		FAB_PG_REQ_HYS,
		FAB_UG_REQ,

		FET_OFF,
		FET_ON,
		FET_OFF_ACK,
		FET_ON_ACK,

		SIP_SAVE_REQ,
		SIP_SAVE_ACK,
		SIP_RESTORE_REQ,
		SIP_RESTORE_ACK,

		SIP_PG_REQ, //PGCB
		SIP_UG_REQ, //PGCB
		FAB_IDLE, //PGCB
		FAB_IDLE_EXIT,//PGCB
		FAB_PG_ACK, //PGCB
		FAB_PG_ACK_DSD,//PGCB
		FAB_PG_NACK,//PGCB
		FAB_PG_NACK_DSD,	//PGCB

		PMC_SIP_WAKE_ALL,
		DEASSERT_PMC_SIP_WAKE_ALL,
		SIP_PG_FLOW,
		SIP_UG_FLOW,
				
		SIP_INACC_PG,
		SIP_INACC_POK,
	
		FAB_PG_FLOW,
		FAB_UG_FLOW,
		PMC_FAB_UG_ALL,

		SET_FET_ON_MODE,
		RESET_FET_ON_MODE,

		AON_SIDE_POK_ASD,

		PRIM_POK_ASD,
		SIDE_POK_ASD,
		PRIM_POK_DSD,
		SIDE_POK_DSD,
	
		PRIM_RST_DSD,
		SIDE_RST_DSD,
		PRIM_RST_ASD,
		SIDE_RST_ASD,

		VNN_ACK_ASD,
		VNN_ACK_DSD,
		VNN_REQ_ASD,
		VNN_REQ_DSD,

		FDFX_BYPASS_ASD,
		FDFX_BYPASS_DSD,
		FDFX_OVR_ASD,
		FDFX_OVR_DSD,

		D3_ASD,
		D3_DSD,
		D0I3_ASD,
		D0I3_DSD

		} Event_e;

/*	typedef enum {
		SIP_IN_ACC,
		WAIT_FOR_SIP_UG_REQ,
		WAIT_FOR_PMC_WAKE_DE,
		WAIT_FOR_SIP_FET_EN,
		WAIT_FOR_SIP_FET_EN_ACK,
		WAIT_FOR_SIP_UG_ACK,
		//RESTORE
		WAIT_FOR_SIP_RESTORE,
		WAIT_FOR_SIP_RESTORE_DSD,
		//RESTORE
		SIP_ON,
		WAIT_FOR_SIP_PG_REQ,
		WAIT_FOR_SIP_PG_ACK,
		SIP_ACC,
		WAIT_FOR_SIP_POK,
		WAIT_FOR_SIP_AON_POK_ASD,
		WAIT_FOR_SIP_POK_DSTD,
		WAIT_FOR_SIP_PG_REQ_INACC,
		WAIT_FOR_SIP_PG_ACK_INACC
		

	} SIPState;
*/
	typedef enum {
		FAB_ON,
		WAIT_FOR_FAB_HYS,
		WAIT_FOR_FAB_ACK_NACK_1,
		WAIT_FOR_FAB_NACK_1,
		WAIT_FOR_FAB_REQ_0_NACK,
		WAIT_FOR_FAB_NACK_0,
		FAB_PG,
		WAIT_FOR_FAB_FET_EN,
		WAIT_FOR_FAB_FET_EN_ACK,		
		WAIT_FOR_FAB_REQ_0_ACK,
		WAIT_FOR_FAB_ACK_0

	} FabricState;


	typedef enum {

		//SIP state
		PWRON,
		PG_REQ,
		PG_HS,
		ACPOF,
		INAPN,
		UGWK_W,
		PGHSI,
		INAPF,
		UGWAK,
		UGFET,
		UGFEA,
		UGHSI,
		UG_REQ,
		UG_HS,
		POKAS,
		POKRS,
		RESTO,

		//fabric
		IDHYS,
		ACKID,
		PWRGT,
		IDEXI,
		ACKEX,
		NACK0,
		REQ_1,
		NACK1,

		//SIP
		INACCESSIBLE_PON,
		INACCESSIBLE_POFF,
		ACCESSIBLE_POFF,
		ACCESSIBLE_PON

		} MonitorState;

	typedef enum {
		SIG,
		MSG,
		SIP,
		FAB,
		FET,
		POK
		} Cycle;

   typedef enum {
		POWER_GATED,
		POWER_UNGATED,
		POWER_UNGATED_POK0
	   } InitialState;

	typedef enum {
		CSME,
		HOST,
		DUAL
	} SIPType;

	typedef enum {
		PHASE_1,
		PHASE_2,
		PHASE_3
	} Phase;
endclass: PowerGating


