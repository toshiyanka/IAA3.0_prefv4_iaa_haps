  `include "hqm_pcie_base_test.sv"
  `include "hqm_pcie_cfg_test.sv"
  `include "hqm_pcie_cfg_error_test.sv"
  `include "hqm_pcie_d3_err_chk_test.sv"
  `include "hqm_pcie_mem_error_test.sv"
  `include "hqm_pcie_error_pollution_test.sv"
  `include "hqm_pcie_cpl_error_test.sv"
  `include "hqm_pcie_tag_test.sv"
  `include "hqm_pcie_mem_test.sv"
  `include "hqm_pcie_hcw_enqueue_test.sv"
  `include "hqm_pcie_unsupported_req_test.sv"
  `include "hqm_pcie_flr_test.sv"
  `include "hqm_pcie_cold_rst_test.sv"
  `include "hqm_pcie_mem_zero_length_read_test.sv"
  `include "hqm_pcie_bypass_np_req_test.sv"
  `include "hqm_pcie_reg_reset_val_test.sv"
  `include "hqm_pcie_flr_with_txns.sv"
  `include "hqm_tlp_rsvd_tgl_test.sv"
  `include "hqm_pcie_cfg_header_check_test.sv"
  `include "hqm_err_report_dis_test.sv"
  `include "hqm_pcie_b2b_single_err_test.sv"
  `include "hqm_tlp_length_test.sv"
  `include "hqm_tlp_fbe_lbe_test.sv"
  `include "hqm_cmd_test.sv"
  `include "hqm_pcie_bar_size_check_test.sv"
  `include "hqm_pasid_variation_test.sv"
  //`include "hqm_pcie_rsvd_type_test.sv"
