module ctech_lib_tieoff_0 (out);
   output logic out;
   d04rid10nnz00 ctech_lib_dcszo (.o(out));
endmodule
