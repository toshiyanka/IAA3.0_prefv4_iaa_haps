`ifndef __VISA_IT__
`ifndef INTEL_GLOBAL_VISA_DISABLE

(* inserted_by="VISA IT" *) logic [162:0] visaPrbsFrom_hqm_core_visa_block;



`endif // INTEL_GLOBAL_VISA_DISABLE
`endif // __VISA_IT__
