case (Node)
   'd0 : begin
            Tap_Info_Int.Next_Tap[0] = NOTAP;
        end
endcase


